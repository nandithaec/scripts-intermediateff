module c499 (
	N1, 
	N5, 
	N9, 
	N13, 
	N17, 
	N21, 
	N25, 
	N29, 
	N33, 
	N37, 
	N41, 
	N45, 
	N49, 
	N53, 
	N57, 
	N61, 
	N65, 
	N69, 
	N73, 
	N77, 
	N81, 
	N85, 
	N89, 
	N93, 
	N97, 
	N101, 
	N105, 
	N109, 
	N113, 
	N117, 
	N121, 
	N125, 
	N129, 
	N130, 
	N131, 
	N132, 
	N133, 
	N134, 
	N135, 
	N136, 
	N137, 
	N724, 
	N725, 
	N726, 
	N727, 
	N728, 
	N729, 
	N730, 
	N731, 
	N732, 
	N733, 
	N734, 
	N735, 
	N736, 
	N737, 
	N738, 
	N739, 
	N740, 
	N741, 
	N742, 
	N743, 
	N744, 
	N745, 
	N746, 
	N747, 
	N748, 
	N749, 
	N750, 
	N751, 
	N752, 
	N753, 
	N754, 
	N755);
   input N1;
   input N5;
   input N9;
   input N13;
   input N17;
   input N21;
   input N25;
   input N29;
   input N33;
   input N37;
   input N41;
   input N45;
   input N49;
   input N53;
   input N57;
   input N61;
   input N65;
   input N69;
   input N73;
   input N77;
   input N81;
   input N85;
   input N89;
   input N93;
   input N97;
   input N101;
   input N105;
   input N109;
   input N113;
   input N117;
   input N121;
   input N125;
   input N129;
   input N130;
   input N131;
   input N132;
   input N133;
   input N134;
   input N135;
   input N136;
   input N137;
   output N724;
   output N725;
   output N726;
   output N727;
   output N728;
   output N729;
   output N730;
   output N731;
   output N732;
   output N733;
   output N734;
   output N735;
   output N736;
   output N737;
   output N738;
   output N739;
   output N740;
   output N741;
   output N742;
   output N743;
   output N744;
   output N745;
   output N746;
   output N747;
   output N748;
   output N749;
   output N750;
   output N751;
   output N752;
   output N753;
   output N754;
   output N755;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;

   INVX2 U1 (.Y(n1), 
	.A(n46));
   INVX2 U2 (.Y(n2), 
	.A(n28));
   INVX2 U3 (.Y(n3), 
	.A(n39));
   INVX2 U4 (.Y(n4), 
	.A(n64));
   INVX2 U5 (.Y(n5), 
	.A(n35));
   INVX2 U6 (.Y(n6), 
	.A(n45));
   INVX2 U7 (.Y(n7), 
	.A(n30));
   INVX2 U8 (.Y(n8), 
	.A(n62));
   INVX2 U9 (.Y(n9), 
	.A(n70));
   INVX2 U10 (.Y(n10), 
	.A(n67));
   INVX2 U11 (.Y(n11), 
	.A(n32));
   INVX2 U12 (.Y(n12), 
	.A(n37));
   INVX2 U13 (.Y(n13), 
	.A(N49));
   INVX2 U14 (.Y(n14), 
	.A(N65));
   INVX2 U15 (.Y(n15), 
	.A(N117));
   XNOR2X1 U16 (.Y(N755), 
	.B(n16), 
	.A(N125));
   NAND2X1 U17 (.Y(n16), 
	.B(n11), 
	.A(n17));
   XNOR2X1 U18 (.Y(N754), 
	.B(n18), 
	.A(N121));
   NAND2X1 U19 (.Y(n18), 
	.B(n5), 
	.A(n17));
   XOR2X1 U20 (.Y(N753), 
	.B(n19), 
	.A(n15));
   NAND2X1 U21 (.Y(n19), 
	.B(n12), 
	.A(n17));
   XNOR2X1 U22 (.Y(N752), 
	.B(n20), 
	.A(N113));
   NAND2X1 U23 (.Y(n20), 
	.B(n3), 
	.A(n17));
   AND2X1 U24 (.Y(n17), 
	.B(n21), 
	.A(n2));
   XNOR2X1 U25 (.Y(N751), 
	.B(n22), 
	.A(N109));
   NAND2X1 U26 (.Y(n22), 
	.B(n11), 
	.A(n23));
   XNOR2X1 U27 (.Y(N750), 
	.B(n24), 
	.A(N105));
   NAND2X1 U28 (.Y(n24), 
	.B(n5), 
	.A(n23));
   XNOR2X1 U29 (.Y(N749), 
	.B(n25), 
	.A(N101));
   NAND2X1 U30 (.Y(n25), 
	.B(n12), 
	.A(n23));
   XNOR2X1 U31 (.Y(N748), 
	.B(n26), 
	.A(N97));
   NAND2X1 U32 (.Y(n26), 
	.B(n3), 
	.A(n23));
   AND2X1 U33 (.Y(n23), 
	.B(n2), 
	.A(n27));
   NAND3X1 U34 (.Y(n28), 
	.C(n30), 
	.B(n29), 
	.A(n8));
   XOR2X1 U35 (.Y(N747), 
	.B(n31), 
	.A(N93));
   NOR2X1 U36 (.Y(n31), 
	.B(n33), 
	.A(n32));
   XOR2X1 U37 (.Y(N746), 
	.B(n34), 
	.A(N89));
   NOR2X1 U38 (.Y(n34), 
	.B(n33), 
	.A(n35));
   XOR2X1 U39 (.Y(N745), 
	.B(n36), 
	.A(N85));
   NOR2X1 U40 (.Y(n36), 
	.B(n33), 
	.A(n37));
   XOR2X1 U41 (.Y(N744), 
	.B(n38), 
	.A(N81));
   NOR2X1 U42 (.Y(n38), 
	.B(n33), 
	.A(n39));
   NAND3X1 U43 (.Y(n33), 
	.C(n6), 
	.B(n29), 
	.A(n21));
   XOR2X1 U44 (.Y(N743), 
	.B(n40), 
	.A(N77));
   NOR2X1 U45 (.Y(n40), 
	.B(n41), 
	.A(n32));
   XOR2X1 U46 (.Y(N742), 
	.B(n42), 
	.A(N73));
   NOR2X1 U47 (.Y(n42), 
	.B(n41), 
	.A(n35));
   XOR2X1 U48 (.Y(N741), 
	.B(n43), 
	.A(N69));
   NOR2X1 U49 (.Y(n43), 
	.B(n41), 
	.A(n37));
   XOR2X1 U50 (.Y(N740), 
	.B(n44), 
	.A(N65));
   NOR2X1 U51 (.Y(n44), 
	.B(n41), 
	.A(n39));
   NAND3X1 U52 (.Y(n41), 
	.C(n6), 
	.B(n29), 
	.A(n27));
   OAI21X1 U53 (.Y(n29), 
	.C(n48), 
	.B(n47), 
	.A(n46));
   NAND2X1 U54 (.Y(n48), 
	.B(n49), 
	.A(n39));
   OAI21X1 U55 (.Y(n49), 
	.C(n50), 
	.B(n5), 
	.A(n11));
   OAI21X1 U56 (.Y(n50), 
	.C(n37), 
	.B(n52), 
	.A(n51));
   NAND2X1 U57 (.Y(n47), 
	.B(n32), 
	.A(n35));
   XNOR2X1 U58 (.Y(N739), 
	.B(n53), 
	.A(N61));
   NAND2X1 U59 (.Y(n53), 
	.B(n10), 
	.A(n54));
   XNOR2X1 U60 (.Y(N738), 
	.B(n55), 
	.A(N57));
   NAND2X1 U61 (.Y(n55), 
	.B(n9), 
	.A(n54));
   XNOR2X1 U62 (.Y(N737), 
	.B(n56), 
	.A(N53));
   NAND2X1 U63 (.Y(n56), 
	.B(n8), 
	.A(n54));
   XOR2X1 U64 (.Y(N736), 
	.B(n57), 
	.A(n13));
   NAND2X1 U65 (.Y(n57), 
	.B(n7), 
	.A(n54));
   AND2X1 U66 (.Y(n54), 
	.B(n51), 
	.A(n4));
   XNOR2X1 U67 (.Y(N735), 
	.B(n58), 
	.A(N45));
   NAND2X1 U68 (.Y(n58), 
	.B(n10), 
	.A(n59));
   XNOR2X1 U69 (.Y(N734), 
	.B(n60), 
	.A(N41));
   NAND2X1 U70 (.Y(n60), 
	.B(n9), 
	.A(n59));
   XNOR2X1 U71 (.Y(N733), 
	.B(n61), 
	.A(N37));
   NAND2X1 U72 (.Y(n61), 
	.B(n8), 
	.A(n59));
   XNOR2X1 U73 (.Y(N732), 
	.B(n63), 
	.A(N33));
   NAND2X1 U74 (.Y(n63), 
	.B(n7), 
	.A(n59));
   AND2X1 U75 (.Y(n59), 
	.B(n4), 
	.A(n52));
   NAND3X1 U76 (.Y(n64), 
	.C(n39), 
	.B(n65), 
	.A(n12));
   XOR2X1 U77 (.Y(N731), 
	.B(n66), 
	.A(N29));
   NOR2X1 U78 (.Y(n66), 
	.B(n68), 
	.A(n67));
   XOR2X1 U79 (.Y(N730), 
	.B(n69), 
	.A(N25));
   NOR2X1 U80 (.Y(n69), 
	.B(n68), 
	.A(n70));
   XOR2X1 U81 (.Y(N729), 
	.B(n71), 
	.A(N21));
   NOR2X1 U82 (.Y(n71), 
	.B(n68), 
	.A(n62));
   XOR2X1 U83 (.Y(N728), 
	.B(n72), 
	.A(N17));
   NOR2X1 U84 (.Y(n72), 
	.B(n68), 
	.A(n30));
   NAND3X1 U85 (.Y(n68), 
	.C(n51), 
	.B(n65), 
	.A(n1));
   NOR2X1 U86 (.Y(n51), 
	.B(n32), 
	.A(n5));
   XOR2X1 U87 (.Y(N727), 
	.B(n73), 
	.A(N13));
   NOR2X1 U88 (.Y(n73), 
	.B(n74), 
	.A(n67));
   XOR2X1 U89 (.Y(N726), 
	.B(n75), 
	.A(N9));
   NOR2X1 U90 (.Y(n75), 
	.B(n74), 
	.A(n70));
   XOR2X1 U91 (.Y(N725), 
	.B(n76), 
	.A(N5));
   NOR2X1 U92 (.Y(n76), 
	.B(n74), 
	.A(n62));
   XOR2X1 U93 (.Y(N724), 
	.B(n77), 
	.A(N1));
   NOR2X1 U94 (.Y(n77), 
	.B(n74), 
	.A(n30));
   NAND3X1 U95 (.Y(n74), 
	.C(n52), 
	.B(n65), 
	.A(n1));
   NOR2X1 U96 (.Y(n52), 
	.B(n35), 
	.A(n11));
   XOR2X1 U97 (.Y(n35), 
	.B(n79), 
	.A(n78));
   XOR2X1 U98 (.Y(n79), 
	.B(n81), 
	.A(n80));
   XOR2X1 U99 (.Y(n81), 
	.B(N105), 
	.A(N121));
   XOR2X1 U100 (.Y(n80), 
	.B(N73), 
	.A(N89));
   XOR2X1 U101 (.Y(n78), 
	.B(n83), 
	.A(n82));
   XOR2X1 U102 (.Y(n82), 
	.B(n85), 
	.A(n84));
   NAND2X1 U103 (.Y(n84), 
	.B(N137), 
	.A(N135));
   XOR2X1 U104 (.Y(n32), 
	.B(n87), 
	.A(n86));
   XOR2X1 U105 (.Y(n87), 
	.B(n89), 
	.A(n88));
   XOR2X1 U106 (.Y(n89), 
	.B(N109), 
	.A(N125));
   XOR2X1 U107 (.Y(n88), 
	.B(N77), 
	.A(N93));
   XOR2X1 U108 (.Y(n86), 
	.B(n91), 
	.A(n90));
   XOR2X1 U109 (.Y(n90), 
	.B(n93), 
	.A(n92));
   NAND2X1 U110 (.Y(n92), 
	.B(N137), 
	.A(N136));
   OAI21X1 U111 (.Y(n65), 
	.C(n95), 
	.B(n94), 
	.A(n45));
   NAND2X1 U112 (.Y(n95), 
	.B(n96), 
	.A(n30));
   OAI21X1 U113 (.Y(n96), 
	.C(n97), 
	.B(n10), 
	.A(n9));
   OAI21X1 U114 (.Y(n97), 
	.C(n62), 
	.B(n27), 
	.A(n21));
   NOR2X1 U115 (.Y(n27), 
	.B(n70), 
	.A(n10));
   NOR2X1 U116 (.Y(n21), 
	.B(n67), 
	.A(n9));
   NAND2X1 U117 (.Y(n94), 
	.B(n67), 
	.A(n70));
   XOR2X1 U118 (.Y(n67), 
	.B(n99), 
	.A(n98));
   XOR2X1 U119 (.Y(n99), 
	.B(n101), 
	.A(n100));
   XOR2X1 U120 (.Y(n101), 
	.B(N13), 
	.A(N29));
   XOR2X1 U121 (.Y(n100), 
	.B(N45), 
	.A(N61));
   XOR2X1 U122 (.Y(n98), 
	.B(n103), 
	.A(n102));
   XOR2X1 U123 (.Y(n102), 
	.B(n105), 
	.A(n104));
   NAND2X1 U124 (.Y(n104), 
	.B(N137), 
	.A(N132));
   XOR2X1 U125 (.Y(n70), 
	.B(n107), 
	.A(n106));
   XOR2X1 U126 (.Y(n107), 
	.B(n109), 
	.A(n108));
   XOR2X1 U127 (.Y(n109), 
	.B(N25), 
	.A(N41));
   XOR2X1 U128 (.Y(n108), 
	.B(N57), 
	.A(N9));
   XOR2X1 U129 (.Y(n106), 
	.B(n111), 
	.A(n110));
   XOR2X1 U130 (.Y(n110), 
	.B(n113), 
	.A(n112));
   NAND2X1 U131 (.Y(n112), 
	.B(N137), 
	.A(N131));
   NAND2X1 U132 (.Y(n45), 
	.B(n7), 
	.A(n62));
   XOR2X1 U133 (.Y(n62), 
	.B(n115), 
	.A(n114));
   XOR2X1 U134 (.Y(n115), 
	.B(n117), 
	.A(n116));
   XOR2X1 U135 (.Y(n117), 
	.B(N21), 
	.A(N37));
   XOR2X1 U136 (.Y(n116), 
	.B(N5), 
	.A(N53));
   XOR2X1 U137 (.Y(n114), 
	.B(n111), 
	.A(n118));
   XNOR2X1 U138 (.Y(n111), 
	.B(n120), 
	.A(n119));
   XOR2X1 U139 (.Y(n120), 
	.B(N109), 
	.A(N97));
   XNOR2X1 U140 (.Y(n119), 
	.B(N105), 
	.A(N101));
   XOR2X1 U141 (.Y(n118), 
	.B(n103), 
	.A(n121));
   XNOR2X1 U142 (.Y(n103), 
	.B(n123), 
	.A(n122));
   XOR2X1 U143 (.Y(n123), 
	.B(N121), 
	.A(N125));
   XOR2X1 U144 (.Y(n122), 
	.B(n15), 
	.A(N113));
   NAND2X1 U145 (.Y(n121), 
	.B(N137), 
	.A(N130));
   NAND2X1 U146 (.Y(n46), 
	.B(n3), 
	.A(n37));
   XOR2X1 U147 (.Y(n39), 
	.B(n125), 
	.A(n124));
   XOR2X1 U148 (.Y(n125), 
	.B(n127), 
	.A(n126));
   XOR2X1 U149 (.Y(n127), 
	.B(N113), 
	.A(N65));
   XOR2X1 U150 (.Y(n126), 
	.B(N81), 
	.A(N97));
   XOR2X1 U151 (.Y(n124), 
	.B(n85), 
	.A(n128));
   XNOR2X1 U152 (.Y(n85), 
	.B(n130), 
	.A(n129));
   XOR2X1 U153 (.Y(n130), 
	.B(N5), 
	.A(N9));
   XNOR2X1 U154 (.Y(n129), 
	.B(N13), 
	.A(N1));
   XOR2X1 U155 (.Y(n128), 
	.B(n93), 
	.A(n131));
   XNOR2X1 U156 (.Y(n93), 
	.B(n133), 
	.A(n132));
   XOR2X1 U157 (.Y(n133), 
	.B(N25), 
	.A(N29));
   XNOR2X1 U158 (.Y(n132), 
	.B(N21), 
	.A(N17));
   NAND2X1 U159 (.Y(n131), 
	.B(N137), 
	.A(N133));
   XOR2X1 U160 (.Y(n37), 
	.B(n135), 
	.A(n134));
   XOR2X1 U161 (.Y(n135), 
	.B(n137), 
	.A(n136));
   XOR2X1 U162 (.Y(n137), 
	.B(N101), 
	.A(N117));
   XOR2X1 U163 (.Y(n136), 
	.B(N69), 
	.A(N85));
   XOR2X1 U164 (.Y(n134), 
	.B(n83), 
	.A(n138));
   XNOR2X1 U165 (.Y(n83), 
	.B(n140), 
	.A(n139));
   XOR2X1 U166 (.Y(n140), 
	.B(N41), 
	.A(N45));
   XNOR2X1 U167 (.Y(n139), 
	.B(N37), 
	.A(N33));
   XOR2X1 U168 (.Y(n138), 
	.B(n91), 
	.A(n141));
   XNOR2X1 U169 (.Y(n91), 
	.B(n143), 
	.A(n142));
   XOR2X1 U170 (.Y(n143), 
	.B(N57), 
	.A(N61));
   XOR2X1 U171 (.Y(n142), 
	.B(N53), 
	.A(n13));
   NAND2X1 U172 (.Y(n141), 
	.B(N134), 
	.A(N137));
   XOR2X1 U173 (.Y(n30), 
	.B(n145), 
	.A(n144));
   XOR2X1 U174 (.Y(n145), 
	.B(n147), 
	.A(n146));
   XOR2X1 U175 (.Y(n147), 
	.B(N1), 
	.A(N17));
   XOR2X1 U176 (.Y(n146), 
	.B(N33), 
	.A(N49));
   XOR2X1 U177 (.Y(n144), 
	.B(n113), 
	.A(n148));
   XNOR2X1 U178 (.Y(n113), 
	.B(n150), 
	.A(n149));
   XOR2X1 U179 (.Y(n150), 
	.B(N73), 
	.A(N77));
   XOR2X1 U180 (.Y(n149), 
	.B(N69), 
	.A(n14));
   XOR2X1 U181 (.Y(n148), 
	.B(n105), 
	.A(n151));
   XNOR2X1 U182 (.Y(n105), 
	.B(n153), 
	.A(n152));
   XOR2X1 U183 (.Y(n153), 
	.B(N89), 
	.A(N93));
   XNOR2X1 U184 (.Y(n152), 
	.B(N85), 
	.A(N81));
   NAND2X1 U185 (.Y(n151), 
	.B(N137), 
	.A(N129));
endmodule

module dff_104 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_103 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_102 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_101 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_100 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_99 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_98 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_97 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_96 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_95 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_94 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_93 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_92 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_91 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_90 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_89 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_88 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_87 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_86 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_85 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_84 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_83 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_82 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_81 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_80 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_79 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_78 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_77 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_76 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_75 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_74 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_73 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_72 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_71 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_70 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_69 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_68 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_67 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_66 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_65 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_64 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_63 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_62 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_61 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_60 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_59 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_58 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_57 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_56 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_55 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_54 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_53 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_52 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_51 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_50 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_49 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_48 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_47 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_46 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_45 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_44 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_43 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_42 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_41 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_40 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_39 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_38 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_37 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_36 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_35 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_34 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_33 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_32 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_31 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_30 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_29 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_28 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_27 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_26 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_25 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_24 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_23 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_22 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_21 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_20 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_19 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_18 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_17 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_16 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_15 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_14 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_13 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_12 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_11 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_10 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_9 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_8 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_7 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_6 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_5 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_4 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_3 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_2 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_1 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module dff_0 (
	q, 
	d, 
	clk);
   output q;
   input d;
   input clk;

   DFFPOSX1 q_reg (.Q(q), 
	.D(d), 
	.CLK(clk));
endmodule

module c499_clk_opFF (
	clk, 
	N1, 
	N5, 
	N9, 
	N13, 
	N17, 
	N21, 
	N25, 
	N29, 
	N33, 
	N37, 
	N41, 
	N45, 
	N49, 
	N53, 
	N57, 
	N61, 
	N65, 
	N69, 
	N73, 
	N77, 
	N81, 
	N85, 
	N89, 
	N93, 
	N97, 
	N101, 
	N105, 
	N109, 
	N113, 
	N117, 
	N121, 
	N125, 
	N129, 
	N130, 
	N131, 
	N132, 
	N133, 
	N134, 
	N135, 
	N136, 
	N137, 
	Qout_N724, 
	Qout_N725, 
	Qout_N726, 
	Qout_N727, 
	Qout_N728, 
	Qout_N729, 
	Qout_N730, 
	Qout_N731, 
	Qout_N732, 
	Qout_N733, 
	Qout_N734, 
	Qout_N735, 
	Qout_N736, 
	Qout_N737, 
	Qout_N738, 
	Qout_N739, 
	Qout_N740, 
	Qout_N741, 
	Qout_N742, 
	Qout_N743, 
	Qout_N744, 
	Qout_N745, 
	Qout_N746, 
	Qout_N747, 
	Qout_N748, 
	Qout_N749, 
	Qout_N750, 
	Qout_N751, 
	Qout_N752, 
	Qout_N753, 
	Qout_N754, 
	Qout_N755);
   input clk;
   input N1;
   input N5;
   input N9;
   input N13;
   input N17;
   input N21;
   input N25;
   input N29;
   input N33;
   input N37;
   input N41;
   input N45;
   input N49;
   input N53;
   input N57;
   input N61;
   input N65;
   input N69;
   input N73;
   input N77;
   input N81;
   input N85;
   input N89;
   input N93;
   input N97;
   input N101;
   input N105;
   input N109;
   input N113;
   input N117;
   input N121;
   input N125;
   input N129;
   input N130;
   input N131;
   input N132;
   input N133;
   input N134;
   input N135;
   input N136;
   input N137;
   output Qout_N724;
   output Qout_N725;
   output Qout_N726;
   output Qout_N727;
   output Qout_N728;
   output Qout_N729;
   output Qout_N730;
   output Qout_N731;
   output Qout_N732;
   output Qout_N733;
   output Qout_N734;
   output Qout_N735;
   output Qout_N736;
   output Qout_N737;
   output Qout_N738;
   output Qout_N739;
   output Qout_N740;
   output Qout_N741;
   output Qout_N742;
   output Qout_N743;
   output Qout_N744;
   output Qout_N745;
   output Qout_N746;
   output Qout_N747;
   output Qout_N748;
   output Qout_N749;
   output Qout_N750;
   output Qout_N751;
   output Qout_N752;
   output Qout_N753;
   output Qout_N754;
   output Qout_N755;

   // Internal wires
   wire clk__L2_N2;
   wire clk__L2_N1;
   wire clk__L2_N0;
   wire clk__L1_N0;
   wire IN_N1;
   wire IN_N5;
   wire IN_N9;
   wire IN_N13;
   wire IN_N17;
   wire IN_N21;
   wire IN_N25;
   wire IN_N29;
   wire IN_N33;
   wire IN_N37;
   wire IN_N41;
   wire IN_N45;
   wire IN_N49;
   wire IN_N53;
   wire IN_N57;
   wire IN_N61;
   wire IN_N65;
   wire IN_N69;
   wire IN_N73;
   wire IN_N77;
   wire IN_N81;
   wire IN_N85;
   wire IN_N89;
   wire IN_N93;
   wire IN_N97;
   wire IN_N101;
   wire IN_N105;
   wire IN_N109;
   wire IN_N113;
   wire IN_N117;
   wire IN_N121;
   wire IN_N125;
   wire IN_N129;
   wire IN_N130;
   wire IN_N131;
   wire IN_N132;
   wire IN_N133;
   wire IN_N134;
   wire IN_N135;
   wire IN_N136;
   wire IN_N137;
   wire N724;
   wire N725;
   wire N726;
   wire N727;
   wire N728;
   wire N729;
   wire N730;
   wire N731;
   wire N732;
   wire N733;
   wire N734;
   wire N735;
   wire N736;
   wire N737;
   wire N738;
   wire N739;
   wire N740;
   wire N741;
   wire N742;
   wire N743;
   wire N744;
   wire N745;
   wire N746;
   wire N747;
   wire N748;
   wire N749;
   wire N750;
   wire N751;
   wire N752;
   wire N753;
   wire N754;
   wire N755;
   wire Q_N724;
   wire Q_N725;
   wire Q_N726;
   wire Q_N727;
   wire Q_N728;
   wire Q_N729;
   wire Q_N730;
   wire Q_N731;
   wire Q_N732;
   wire Q_N733;
   wire Q_N734;
   wire Q_N735;
   wire Q_N736;
   wire Q_N737;
   wire Q_N738;
   wire Q_N739;
   wire Q_N740;
   wire Q_N741;
   wire Q_N742;
   wire Q_N743;
   wire Q_N744;
   wire Q_N745;
   wire Q_N746;
   wire Q_N747;
   wire Q_N748;
   wire Q_N749;
   wire Q_N750;
   wire Q_N751;
   wire Q_N752;
   wire Q_N753;
   wire Q_N754;
   wire Q_N755;

   INVX8 clk__L2_I2 (.Y(clk__L2_N2), 
	.A(clk__L1_N0));
   INVX8 clk__L2_I1 (.Y(clk__L2_N1), 
	.A(clk__L1_N0));
   INVX8 clk__L2_I0 (.Y(clk__L2_N0), 
	.A(clk__L1_N0));
   INVX8 clk__L1_I0 (.Y(clk__L1_N0), 
	.A(clk));
   c499 c0 (.N1(IN_N1), 
	.N5(IN_N5), 
	.N9(IN_N9), 
	.N13(IN_N13), 
	.N17(IN_N17), 
	.N21(IN_N21), 
	.N25(IN_N25), 
	.N29(IN_N29), 
	.N33(IN_N33), 
	.N37(IN_N37), 
	.N41(IN_N41), 
	.N45(IN_N45), 
	.N49(IN_N49), 
	.N53(IN_N53), 
	.N57(IN_N57), 
	.N61(IN_N61), 
	.N65(IN_N65), 
	.N69(IN_N69), 
	.N73(IN_N73), 
	.N77(IN_N77), 
	.N81(IN_N81), 
	.N85(IN_N85), 
	.N89(IN_N89), 
	.N93(IN_N93), 
	.N97(IN_N97), 
	.N101(IN_N101), 
	.N105(IN_N105), 
	.N109(IN_N109), 
	.N113(IN_N113), 
	.N117(IN_N117), 
	.N121(IN_N121), 
	.N125(IN_N125), 
	.N129(IN_N129), 
	.N130(IN_N130), 
	.N131(IN_N131), 
	.N132(IN_N132), 
	.N133(IN_N133), 
	.N134(IN_N134), 
	.N135(IN_N135), 
	.N136(IN_N136), 
	.N137(IN_N137), 
	.N724(N724), 
	.N725(N725), 
	.N726(N726), 
	.N727(N727), 
	.N728(N728), 
	.N729(N729), 
	.N730(N730), 
	.N731(N731), 
	.N732(N732), 
	.N733(N733), 
	.N734(N734), 
	.N735(N735), 
	.N736(N736), 
	.N737(N737), 
	.N738(N738), 
	.N739(N739), 
	.N740(N740), 
	.N741(N741), 
	.N742(N742), 
	.N743(N743), 
	.N744(N744), 
	.N745(N745), 
	.N746(N746), 
	.N747(N747), 
	.N748(N748), 
	.N749(N749), 
	.N750(N750), 
	.N751(N751), 
	.N752(N752), 
	.N753(N753), 
	.N754(N754), 
	.N755(N755));
   dff_104 iDFF_1 (.q(IN_N1), 
	.d(N1), 
	.clk(clk__L2_N2));
   dff_103 iDFF_2 (.q(IN_N5), 
	.d(N5), 
	.clk(clk__L2_N2));
   dff_102 iDFF_3 (.q(IN_N9), 
	.d(N9), 
	.clk(clk__L2_N2));
   dff_101 iDFF_4 (.q(IN_N13), 
	.d(N13), 
	.clk(clk__L2_N2));
   dff_100 iDFF_5 (.q(IN_N17), 
	.d(N17), 
	.clk(clk__L2_N1));
   dff_99 iDFF_6 (.q(IN_N21), 
	.d(N21), 
	.clk(clk__L2_N1));
   dff_98 iDFF_7 (.q(IN_N25), 
	.d(N25), 
	.clk(clk__L2_N2));
   dff_97 iDFF_8 (.q(IN_N29), 
	.d(N29), 
	.clk(clk__L2_N2));
   dff_96 iDFF_9 (.q(IN_N33), 
	.d(N33), 
	.clk(clk__L2_N1));
   dff_95 iDFF_10 (.q(IN_N37), 
	.d(N37), 
	.clk(clk__L2_N1));
   dff_94 iDFF_11 (.q(IN_N41), 
	.d(N41), 
	.clk(clk__L2_N2));
   dff_93 iDFF_12 (.q(IN_N45), 
	.d(N45), 
	.clk(clk__L2_N2));
   dff_92 iDFF_13 (.q(IN_N49), 
	.d(N49), 
	.clk(clk__L2_N1));
   dff_91 iDFF_14 (.q(IN_N53), 
	.d(N53), 
	.clk(clk__L2_N2));
   dff_90 iDFF_15 (.q(IN_N57), 
	.d(N57), 
	.clk(clk__L2_N2));
   dff_89 iDFF_16 (.q(IN_N61), 
	.d(N61), 
	.clk(clk__L2_N2));
   dff_88 iDFF_17 (.q(IN_N65), 
	.d(N65), 
	.clk(clk__L2_N0));
   dff_87 iDFF_18 (.q(IN_N69), 
	.d(N69), 
	.clk(clk__L2_N0));
   dff_86 iDFF_19 (.q(IN_N73), 
	.d(N73), 
	.clk(clk__L2_N0));
   dff_85 iDFF_20 (.q(IN_N77), 
	.d(N77), 
	.clk(clk__L2_N1));
   dff_84 iDFF_21 (.q(IN_N81), 
	.d(N81), 
	.clk(clk__L2_N0));
   dff_83 iDFF_22 (.q(IN_N85), 
	.d(N85), 
	.clk(clk__L2_N0));
   dff_82 iDFF_23 (.q(IN_N89), 
	.d(N89), 
	.clk(clk__L2_N1));
   dff_81 iDFF_24 (.q(IN_N93), 
	.d(N93), 
	.clk(clk__L2_N1));
   dff_80 iDFF_25 (.q(IN_N97), 
	.d(N97), 
	.clk(clk__L2_N0));
   dff_79 iDFF_26 (.q(IN_N101), 
	.d(N101), 
	.clk(clk__L2_N0));
   dff_78 iDFF_27 (.q(IN_N105), 
	.d(N105), 
	.clk(clk__L2_N0));
   dff_77 iDFF_28 (.q(IN_N109), 
	.d(N109), 
	.clk(clk__L2_N0));
   dff_76 iDFF_29 (.q(IN_N113), 
	.d(N113), 
	.clk(clk__L2_N0));
   dff_75 iDFF_30 (.q(IN_N117), 
	.d(N117), 
	.clk(clk__L2_N0));
   dff_74 iDFF_31 (.q(IN_N121), 
	.d(N121), 
	.clk(clk__L2_N1));
   dff_73 iDFF_32 (.q(IN_N125), 
	.d(N125), 
	.clk(clk__L2_N1));
   dff_72 iDFF_33 (.q(IN_N129), 
	.d(N129), 
	.clk(clk__L2_N1));
   dff_71 iDFF_34 (.q(IN_N130), 
	.d(N130), 
	.clk(clk__L2_N1));
   dff_70 iDFF_35 (.q(IN_N131), 
	.d(N131), 
	.clk(clk__L2_N1));
   dff_69 iDFF_36 (.q(IN_N132), 
	.d(N132), 
	.clk(clk__L2_N1));
   dff_68 iDFF_37 (.q(IN_N133), 
	.d(N133), 
	.clk(clk__L2_N1));
   dff_67 iDFF_38 (.q(IN_N134), 
	.d(N134), 
	.clk(clk__L2_N1));
   dff_66 iDFF_39 (.q(IN_N135), 
	.d(N135), 
	.clk(clk__L2_N0));
   dff_65 iDFF_40 (.q(IN_N136), 
	.d(N136), 
	.clk(clk__L2_N1));
   dff_64 iDFF_41 (.q(IN_N137), 
	.d(N137), 
	.clk(clk__L2_N1));
   dff_63 DFF_1 (.q(Q_N724), 
	.d(N724), 
	.clk(clk__L2_N2));
   dff_62 DFF_2 (.q(Q_N725), 
	.d(N725), 
	.clk(clk__L2_N2));
   dff_61 DFF_3 (.q(Q_N726), 
	.d(N726), 
	.clk(clk__L2_N2));
   dff_60 DFF_4 (.q(Q_N727), 
	.d(N727), 
	.clk(clk__L2_N2));
   dff_59 DFF_5 (.q(Q_N728), 
	.d(N728), 
	.clk(clk__L2_N2));
   dff_58 DFF_6 (.q(Q_N729), 
	.d(N729), 
	.clk(clk__L2_N1));
   dff_57 DFF_7 (.q(Q_N730), 
	.d(N730), 
	.clk(clk__L2_N2));
   dff_56 DFF_8 (.q(Q_N731), 
	.d(N731), 
	.clk(clk__L2_N2));
   dff_55 DFF_9 (.q(Q_N732), 
	.d(N732), 
	.clk(clk__L2_N1));
   dff_54 DFF_10 (.q(Q_N733), 
	.d(N733), 
	.clk(clk__L2_N1));
   dff_53 DFF_11 (.q(Q_N734), 
	.d(N734), 
	.clk(clk__L2_N2));
   dff_52 DFF_12 (.q(Q_N735), 
	.d(N735), 
	.clk(clk__L2_N2));
   dff_51 DFF_13 (.q(Q_N736), 
	.d(N736), 
	.clk(clk__L2_N1));
   dff_50 DFF_14 (.q(Q_N737), 
	.d(N737), 
	.clk(clk__L2_N2));
   dff_49 DFF_15 (.q(Q_N738), 
	.d(N738), 
	.clk(clk__L2_N2));
   dff_48 DFF_16 (.q(Q_N739), 
	.d(N739), 
	.clk(clk__L2_N2));
   dff_47 DFF_17 (.q(Q_N740), 
	.d(N740), 
	.clk(clk__L2_N0));
   dff_46 DFF_18 (.q(Q_N741), 
	.d(N741), 
	.clk(clk__L2_N0));
   dff_45 DFF_19 (.q(Q_N742), 
	.d(N742), 
	.clk(clk__L2_N0));
   dff_44 DFF_20 (.q(Q_N743), 
	.d(N743), 
	.clk(clk__L2_N1));
   dff_43 DFF_21 (.q(Q_N744), 
	.d(N744), 
	.clk(clk__L2_N0));
   dff_42 DFF_22 (.q(Q_N745), 
	.d(N745), 
	.clk(clk__L2_N0));
   dff_41 DFF_23 (.q(Q_N746), 
	.d(N746), 
	.clk(clk__L2_N0));
   dff_40 DFF_24 (.q(Q_N747), 
	.d(N747), 
	.clk(clk__L2_N1));
   dff_39 DFF_25 (.q(Q_N748), 
	.d(N748), 
	.clk(clk__L2_N0));
   dff_38 DFF_26 (.q(Q_N749), 
	.d(N749), 
	.clk(clk__L2_N0));
   dff_37 DFF_27 (.q(Q_N750), 
	.d(N750), 
	.clk(clk__L2_N0));
   dff_36 DFF_28 (.q(Q_N751), 
	.d(N751), 
	.clk(clk__L2_N1));
   dff_35 DFF_29 (.q(Q_N752), 
	.d(N752), 
	.clk(clk__L2_N0));
   dff_34 DFF_30 (.q(Q_N753), 
	.d(N753), 
	.clk(clk__L2_N0));
   dff_33 DFF_31 (.q(Q_N754), 
	.d(N754), 
	.clk(clk__L2_N1));
   dff_32 DFF_32 (.q(Q_N755), 
	.d(N755), 
	.clk(clk__L2_N1));
   dff_31 oDFF_1 (.q(Qout_N724), 
	.d(Q_N724), 
	.clk(clk__L2_N2));
   dff_30 oDFF_2 (.q(Qout_N725), 
	.d(Q_N725), 
	.clk(clk__L2_N2));
   dff_29 oDFF_3 (.q(Qout_N726), 
	.d(Q_N726), 
	.clk(clk__L2_N2));
   dff_28 oDFF_4 (.q(Qout_N727), 
	.d(Q_N727), 
	.clk(clk__L2_N2));
   dff_27 oDFF_5 (.q(Qout_N728), 
	.d(Q_N728), 
	.clk(clk__L2_N1));
   dff_26 oDFF_6 (.q(Qout_N729), 
	.d(Q_N729), 
	.clk(clk__L2_N2));
   dff_25 oDFF_7 (.q(Qout_N730), 
	.d(Q_N730), 
	.clk(clk__L2_N2));
   dff_24 oDFF_8 (.q(Qout_N731), 
	.d(Q_N731), 
	.clk(clk__L2_N2));
   dff_23 oDFF_9 (.q(Qout_N732), 
	.d(Q_N732), 
	.clk(clk__L2_N1));
   dff_22 oDFF_10 (.q(Qout_N733), 
	.d(Q_N733), 
	.clk(clk__L2_N1));
   dff_21 oDFF_11 (.q(Qout_N734), 
	.d(Q_N734), 
	.clk(clk__L2_N2));
   dff_20 oDFF_12 (.q(Qout_N735), 
	.d(Q_N735), 
	.clk(clk__L2_N2));
   dff_19 oDFF_13 (.q(Qout_N736), 
	.d(Q_N736), 
	.clk(clk__L2_N1));
   dff_18 oDFF_14 (.q(Qout_N737), 
	.d(Q_N737), 
	.clk(clk__L2_N2));
   dff_17 oDFF_15 (.q(Qout_N738), 
	.d(Q_N738), 
	.clk(clk__L2_N2));
   dff_16 oDFF_16 (.q(Qout_N739), 
	.d(Q_N739), 
	.clk(clk__L2_N2));
   dff_15 oDFF_17 (.q(Qout_N740), 
	.d(Q_N740), 
	.clk(clk__L2_N0));
   dff_14 oDFF_18 (.q(Qout_N741), 
	.d(Q_N741), 
	.clk(clk__L2_N0));
   dff_13 oDFF_19 (.q(Qout_N742), 
	.d(Q_N742), 
	.clk(clk__L2_N0));
   dff_12 oDFF_20 (.q(Qout_N743), 
	.d(Q_N743), 
	.clk(clk__L2_N1));
   dff_11 oDFF_21 (.q(Qout_N744), 
	.d(Q_N744), 
	.clk(clk__L2_N0));
   dff_10 oDFF_22 (.q(Qout_N745), 
	.d(Q_N745), 
	.clk(clk__L2_N0));
   dff_9 oDFF_23 (.q(Qout_N746), 
	.d(Q_N746), 
	.clk(clk__L2_N0));
   dff_8 oDFF_24 (.q(Qout_N747), 
	.d(Q_N747), 
	.clk(clk__L2_N1));
   dff_7 oDFF_25 (.q(Qout_N748), 
	.d(Q_N748), 
	.clk(clk__L2_N0));
   dff_6 oDFF_26 (.q(Qout_N749), 
	.d(Q_N749), 
	.clk(clk__L2_N0));
   dff_5 oDFF_27 (.q(Qout_N750), 
	.d(Q_N750), 
	.clk(clk__L2_N0));
   dff_4 oDFF_28 (.q(Qout_N751), 
	.d(Q_N751), 
	.clk(clk__L2_N1));
   dff_3 oDFF_29 (.q(Qout_N752), 
	.d(Q_N752), 
	.clk(clk__L2_N0));
   dff_2 oDFF_30 (.q(Qout_N753), 
	.d(Q_N753), 
	.clk(clk__L2_N0));
   dff_1 oDFF_31 (.q(Qout_N754), 
	.d(Q_N754), 
	.clk(clk__L2_N0));
   dff_0 oDFF_32 (.q(Qout_N755), 
	.d(Q_N755), 
	.clk(clk__L2_N1));
//************************* CODE APPENDED TO ORIGINAL .v FILE STARTS FROM HERE *************************
integer fileout;
integer clk_count = 0;
integer fileout1;
integer clk_count1 = 0;
initial
begin
fileout= $fopen("./c499_clk_opFF_reference_out/our_reference_out.txt","a+");
fileout1= $fopen("./c499_clk_opFF_reference_out/tool_reference_out.txt","a+");
end
always @(negedge clk)
begin
$fwrite(fileout,"IN_N1 = %b\n", IN_N1);
$fwrite(fileout1,"%b ", IN_N1);
$fwrite(fileout,"IN_N5 = %b\n", IN_N5);
$fwrite(fileout1,"%b ", IN_N5);
$fwrite(fileout,"IN_N9 = %b\n", IN_N9);
$fwrite(fileout1,"%b ", IN_N9);
$fwrite(fileout,"IN_N13 = %b\n", IN_N13);
$fwrite(fileout1,"%b ", IN_N13);
$fwrite(fileout,"IN_N17 = %b\n", IN_N17);
$fwrite(fileout1,"%b ", IN_N17);
$fwrite(fileout,"IN_N21 = %b\n", IN_N21);
$fwrite(fileout1,"%b ", IN_N21);
$fwrite(fileout,"IN_N25 = %b\n", IN_N25);
$fwrite(fileout1,"%b ", IN_N25);
$fwrite(fileout,"IN_N29 = %b\n", IN_N29);
$fwrite(fileout1,"%b ", IN_N29);
$fwrite(fileout,"IN_N33 = %b\n", IN_N33);
$fwrite(fileout1,"%b ", IN_N33);
$fwrite(fileout,"IN_N37 = %b\n", IN_N37);
$fwrite(fileout1,"%b ", IN_N37);
$fwrite(fileout,"IN_N41 = %b\n", IN_N41);
$fwrite(fileout1,"%b ", IN_N41);
$fwrite(fileout,"IN_N45 = %b\n", IN_N45);
$fwrite(fileout1,"%b ", IN_N45);
$fwrite(fileout,"IN_N49 = %b\n", IN_N49);
$fwrite(fileout1,"%b ", IN_N49);
$fwrite(fileout,"IN_N53 = %b\n", IN_N53);
$fwrite(fileout1,"%b ", IN_N53);
$fwrite(fileout,"IN_N57 = %b\n", IN_N57);
$fwrite(fileout1,"%b ", IN_N57);
$fwrite(fileout,"IN_N61 = %b\n", IN_N61);
$fwrite(fileout1,"%b ", IN_N61);
$fwrite(fileout,"IN_N65 = %b\n", IN_N65);
$fwrite(fileout1,"%b ", IN_N65);
$fwrite(fileout,"IN_N69 = %b\n", IN_N69);
$fwrite(fileout1,"%b ", IN_N69);
$fwrite(fileout,"IN_N73 = %b\n", IN_N73);
$fwrite(fileout1,"%b ", IN_N73);
$fwrite(fileout,"IN_N77 = %b\n", IN_N77);
$fwrite(fileout1,"%b ", IN_N77);
$fwrite(fileout,"IN_N81 = %b\n", IN_N81);
$fwrite(fileout1,"%b ", IN_N81);
$fwrite(fileout,"IN_N85 = %b\n", IN_N85);
$fwrite(fileout1,"%b ", IN_N85);
$fwrite(fileout,"IN_N89 = %b\n", IN_N89);
$fwrite(fileout1,"%b ", IN_N89);
$fwrite(fileout,"IN_N93 = %b\n", IN_N93);
$fwrite(fileout1,"%b ", IN_N93);
$fwrite(fileout,"IN_N97 = %b\n", IN_N97);
$fwrite(fileout1,"%b ", IN_N97);
$fwrite(fileout,"IN_N101 = %b\n", IN_N101);
$fwrite(fileout1,"%b ", IN_N101);
$fwrite(fileout,"IN_N105 = %b\n", IN_N105);
$fwrite(fileout1,"%b ", IN_N105);
$fwrite(fileout,"IN_N109 = %b\n", IN_N109);
$fwrite(fileout1,"%b ", IN_N109);
$fwrite(fileout,"IN_N113 = %b\n", IN_N113);
$fwrite(fileout1,"%b ", IN_N113);
$fwrite(fileout,"IN_N117 = %b\n", IN_N117);
$fwrite(fileout1,"%b ", IN_N117);
$fwrite(fileout,"IN_N121 = %b\n", IN_N121);
$fwrite(fileout1,"%b ", IN_N121);
$fwrite(fileout,"IN_N125 = %b\n", IN_N125);
$fwrite(fileout1,"%b ", IN_N125);
$fwrite(fileout,"IN_N129 = %b\n", IN_N129);
$fwrite(fileout1,"%b ", IN_N129);
$fwrite(fileout,"IN_N130 = %b\n", IN_N130);
$fwrite(fileout1,"%b ", IN_N130);
$fwrite(fileout,"IN_N131 = %b\n", IN_N131);
$fwrite(fileout1,"%b ", IN_N131);
$fwrite(fileout,"IN_N132 = %b\n", IN_N132);
$fwrite(fileout1,"%b ", IN_N132);
$fwrite(fileout,"IN_N133 = %b\n", IN_N133);
$fwrite(fileout1,"%b ", IN_N133);
$fwrite(fileout,"IN_N134 = %b\n", IN_N134);
$fwrite(fileout1,"%b ", IN_N134);
$fwrite(fileout,"IN_N135 = %b\n", IN_N135);
$fwrite(fileout1,"%b ", IN_N135);
$fwrite(fileout,"IN_N136 = %b\n", IN_N136);
$fwrite(fileout1,"%b ", IN_N136);
$fwrite(fileout,"IN_N137 = %b\n", IN_N137);
$fwrite(fileout1,"%b ", IN_N137);
$fwrite(fileout,"Q_N724 = %b\n", Q_N724);
$fwrite(fileout1,"%b ", Q_N724);
$fwrite(fileout,"Q_N725 = %b\n", Q_N725);
$fwrite(fileout1,"%b ", Q_N725);
$fwrite(fileout,"Q_N726 = %b\n", Q_N726);
$fwrite(fileout1,"%b ", Q_N726);
$fwrite(fileout,"Q_N727 = %b\n", Q_N727);
$fwrite(fileout1,"%b ", Q_N727);
$fwrite(fileout,"Q_N728 = %b\n", Q_N728);
$fwrite(fileout1,"%b ", Q_N728);
$fwrite(fileout,"Q_N729 = %b\n", Q_N729);
$fwrite(fileout1,"%b ", Q_N729);
$fwrite(fileout,"Q_N730 = %b\n", Q_N730);
$fwrite(fileout1,"%b ", Q_N730);
$fwrite(fileout,"Q_N731 = %b\n", Q_N731);
$fwrite(fileout1,"%b ", Q_N731);
$fwrite(fileout,"Q_N732 = %b\n", Q_N732);
$fwrite(fileout1,"%b ", Q_N732);
$fwrite(fileout,"Q_N733 = %b\n", Q_N733);
$fwrite(fileout1,"%b ", Q_N733);
$fwrite(fileout,"Q_N734 = %b\n", Q_N734);
$fwrite(fileout1,"%b ", Q_N734);
$fwrite(fileout,"Q_N735 = %b\n", Q_N735);
$fwrite(fileout1,"%b ", Q_N735);
$fwrite(fileout,"Q_N736 = %b\n", Q_N736);
$fwrite(fileout1,"%b ", Q_N736);
$fwrite(fileout,"Q_N737 = %b\n", Q_N737);
$fwrite(fileout1,"%b ", Q_N737);
$fwrite(fileout,"Q_N738 = %b\n", Q_N738);
$fwrite(fileout1,"%b ", Q_N738);
$fwrite(fileout,"Q_N739 = %b\n", Q_N739);
$fwrite(fileout1,"%b ", Q_N739);
$fwrite(fileout,"Q_N740 = %b\n", Q_N740);
$fwrite(fileout1,"%b ", Q_N740);
$fwrite(fileout,"Q_N741 = %b\n", Q_N741);
$fwrite(fileout1,"%b ", Q_N741);
$fwrite(fileout,"Q_N742 = %b\n", Q_N742);
$fwrite(fileout1,"%b ", Q_N742);
$fwrite(fileout,"Q_N743 = %b\n", Q_N743);
$fwrite(fileout1,"%b ", Q_N743);
$fwrite(fileout,"Q_N744 = %b\n", Q_N744);
$fwrite(fileout1,"%b ", Q_N744);
$fwrite(fileout,"Q_N745 = %b\n", Q_N745);
$fwrite(fileout1,"%b ", Q_N745);
$fwrite(fileout,"Q_N746 = %b\n", Q_N746);
$fwrite(fileout1,"%b ", Q_N746);
$fwrite(fileout,"Q_N747 = %b\n", Q_N747);
$fwrite(fileout1,"%b ", Q_N747);
$fwrite(fileout,"Q_N748 = %b\n", Q_N748);
$fwrite(fileout1,"%b ", Q_N748);
$fwrite(fileout,"Q_N749 = %b\n", Q_N749);
$fwrite(fileout1,"%b ", Q_N749);
$fwrite(fileout,"Q_N750 = %b\n", Q_N750);
$fwrite(fileout1,"%b ", Q_N750);
$fwrite(fileout,"Q_N751 = %b\n", Q_N751);
$fwrite(fileout1,"%b ", Q_N751);
$fwrite(fileout,"Q_N752 = %b\n", Q_N752);
$fwrite(fileout1,"%b ", Q_N752);
$fwrite(fileout,"Q_N753 = %b\n", Q_N753);
$fwrite(fileout1,"%b ", Q_N753);
$fwrite(fileout,"Q_N754 = %b\n", Q_N754);
$fwrite(fileout1,"%b ", Q_N754);
$fwrite(fileout,"Q_N755 = %b\n", Q_N755);
$fwrite(fileout1,"%b ", Q_N755);
$fwrite(fileout,"Qout_N724 = %b\n", Qout_N724);
$fwrite(fileout1,"%b ", Qout_N724);
$fwrite(fileout,"Qout_N725 = %b\n", Qout_N725);
$fwrite(fileout1,"%b ", Qout_N725);
$fwrite(fileout,"Qout_N726 = %b\n", Qout_N726);
$fwrite(fileout1,"%b ", Qout_N726);
$fwrite(fileout,"Qout_N727 = %b\n", Qout_N727);
$fwrite(fileout1,"%b ", Qout_N727);
$fwrite(fileout,"Qout_N728 = %b\n", Qout_N728);
$fwrite(fileout1,"%b ", Qout_N728);
$fwrite(fileout,"Qout_N729 = %b\n", Qout_N729);
$fwrite(fileout1,"%b ", Qout_N729);
$fwrite(fileout,"Qout_N730 = %b\n", Qout_N730);
$fwrite(fileout1,"%b ", Qout_N730);
$fwrite(fileout,"Qout_N731 = %b\n", Qout_N731);
$fwrite(fileout1,"%b ", Qout_N731);
$fwrite(fileout,"Qout_N732 = %b\n", Qout_N732);
$fwrite(fileout1,"%b ", Qout_N732);
$fwrite(fileout,"Qout_N733 = %b\n", Qout_N733);
$fwrite(fileout1,"%b ", Qout_N733);
$fwrite(fileout,"Qout_N734 = %b\n", Qout_N734);
$fwrite(fileout1,"%b ", Qout_N734);
$fwrite(fileout,"Qout_N735 = %b\n", Qout_N735);
$fwrite(fileout1,"%b ", Qout_N735);
$fwrite(fileout,"Qout_N736 = %b\n", Qout_N736);
$fwrite(fileout1,"%b ", Qout_N736);
$fwrite(fileout,"Qout_N737 = %b\n", Qout_N737);
$fwrite(fileout1,"%b ", Qout_N737);
$fwrite(fileout,"Qout_N738 = %b\n", Qout_N738);
$fwrite(fileout1,"%b ", Qout_N738);
$fwrite(fileout,"Qout_N739 = %b\n", Qout_N739);
$fwrite(fileout1,"%b ", Qout_N739);
$fwrite(fileout,"Qout_N740 = %b\n", Qout_N740);
$fwrite(fileout1,"%b ", Qout_N740);
$fwrite(fileout,"Qout_N741 = %b\n", Qout_N741);
$fwrite(fileout1,"%b ", Qout_N741);
$fwrite(fileout,"Qout_N742 = %b\n", Qout_N742);
$fwrite(fileout1,"%b ", Qout_N742);
$fwrite(fileout,"Qout_N743 = %b\n", Qout_N743);
$fwrite(fileout1,"%b ", Qout_N743);
$fwrite(fileout,"Qout_N744 = %b\n", Qout_N744);
$fwrite(fileout1,"%b ", Qout_N744);
$fwrite(fileout,"Qout_N745 = %b\n", Qout_N745);
$fwrite(fileout1,"%b ", Qout_N745);
$fwrite(fileout,"Qout_N746 = %b\n", Qout_N746);
$fwrite(fileout1,"%b ", Qout_N746);
$fwrite(fileout,"Qout_N747 = %b\n", Qout_N747);
$fwrite(fileout1,"%b ", Qout_N747);
$fwrite(fileout,"Qout_N748 = %b\n", Qout_N748);
$fwrite(fileout1,"%b ", Qout_N748);
$fwrite(fileout,"Qout_N749 = %b\n", Qout_N749);
$fwrite(fileout1,"%b ", Qout_N749);
$fwrite(fileout,"Qout_N750 = %b\n", Qout_N750);
$fwrite(fileout1,"%b ", Qout_N750);
$fwrite(fileout,"Qout_N751 = %b\n", Qout_N751);
$fwrite(fileout1,"%b ", Qout_N751);
$fwrite(fileout,"Qout_N752 = %b\n", Qout_N752);
$fwrite(fileout1,"%b ", Qout_N752);
$fwrite(fileout,"Qout_N753 = %b\n", Qout_N753);
$fwrite(fileout1,"%b ", Qout_N753);
$fwrite(fileout,"Qout_N754 = %b\n", Qout_N754);
$fwrite(fileout1,"%b ", Qout_N754);
$fwrite(fileout,"Qout_N755 = %b\n", Qout_N755);
$fwrite(fileout1,"%b ", Qout_N755);
$fwrite(fileout,"\n");
$fwrite(fileout1,"\n");
$fwrite(fileout,"%d CLOCK CYCLE ENDS   :SIGNAL VALUES AT THIS POINT \n\n",clk_count);
$fwrite(fileout,"***********************************************************************************************************\n\n");
end
always @(posedge clk)
begin
clk_count=clk_count+1;
$fwrite(fileout,"%d CLOCK CYCLE STARTS :SIGNAL VALUES AT THIS POINT \n\n",clk_count);
$fwrite(fileout,"N1 = %b\n", N1);
$fwrite(fileout1,"%b ", N1);
$fwrite(fileout,"N5 = %b\n", N5);
$fwrite(fileout1,"%b ", N5);
$fwrite(fileout,"N9 = %b\n", N9);
$fwrite(fileout1,"%b ", N9);
$fwrite(fileout,"N13 = %b\n", N13);
$fwrite(fileout1,"%b ", N13);
$fwrite(fileout,"N17 = %b\n", N17);
$fwrite(fileout1,"%b ", N17);
$fwrite(fileout,"N21 = %b\n", N21);
$fwrite(fileout1,"%b ", N21);
$fwrite(fileout,"N25 = %b\n", N25);
$fwrite(fileout1,"%b ", N25);
$fwrite(fileout,"N29 = %b\n", N29);
$fwrite(fileout1,"%b ", N29);
$fwrite(fileout,"N33 = %b\n", N33);
$fwrite(fileout1,"%b ", N33);
$fwrite(fileout,"N37 = %b\n", N37);
$fwrite(fileout1,"%b ", N37);
$fwrite(fileout,"N41 = %b\n", N41);
$fwrite(fileout1,"%b ", N41);
$fwrite(fileout,"N45 = %b\n", N45);
$fwrite(fileout1,"%b ", N45);
$fwrite(fileout,"N49 = %b\n", N49);
$fwrite(fileout1,"%b ", N49);
$fwrite(fileout,"N53 = %b\n", N53);
$fwrite(fileout1,"%b ", N53);
$fwrite(fileout,"N57 = %b\n", N57);
$fwrite(fileout1,"%b ", N57);
$fwrite(fileout,"N61 = %b\n", N61);
$fwrite(fileout1,"%b ", N61);
$fwrite(fileout,"N65 = %b\n", N65);
$fwrite(fileout1,"%b ", N65);
$fwrite(fileout,"N69 = %b\n", N69);
$fwrite(fileout1,"%b ", N69);
$fwrite(fileout,"N73 = %b\n", N73);
$fwrite(fileout1,"%b ", N73);
$fwrite(fileout,"N77 = %b\n", N77);
$fwrite(fileout1,"%b ", N77);
$fwrite(fileout,"N81 = %b\n", N81);
$fwrite(fileout1,"%b ", N81);
$fwrite(fileout,"N85 = %b\n", N85);
$fwrite(fileout1,"%b ", N85);
$fwrite(fileout,"N89 = %b\n", N89);
$fwrite(fileout1,"%b ", N89);
$fwrite(fileout,"N93 = %b\n", N93);
$fwrite(fileout1,"%b ", N93);
$fwrite(fileout,"N97 = %b\n", N97);
$fwrite(fileout1,"%b ", N97);
$fwrite(fileout,"N101 = %b\n", N101);
$fwrite(fileout1,"%b ", N101);
$fwrite(fileout,"N105 = %b\n", N105);
$fwrite(fileout1,"%b ", N105);
$fwrite(fileout,"N109 = %b\n", N109);
$fwrite(fileout1,"%b ", N109);
$fwrite(fileout,"N113 = %b\n", N113);
$fwrite(fileout1,"%b ", N113);
$fwrite(fileout,"N117 = %b\n", N117);
$fwrite(fileout1,"%b ", N117);
$fwrite(fileout,"N121 = %b\n", N121);
$fwrite(fileout1,"%b ", N121);
$fwrite(fileout,"N125 = %b\n", N125);
$fwrite(fileout1,"%b ", N125);
$fwrite(fileout,"N129 = %b\n", N129);
$fwrite(fileout1,"%b ", N129);
$fwrite(fileout,"N130 = %b\n", N130);
$fwrite(fileout1,"%b ", N130);
$fwrite(fileout,"N131 = %b\n", N131);
$fwrite(fileout1,"%b ", N131);
$fwrite(fileout,"N132 = %b\n", N132);
$fwrite(fileout1,"%b ", N132);
$fwrite(fileout,"N133 = %b\n", N133);
$fwrite(fileout1,"%b ", N133);
$fwrite(fileout,"N134 = %b\n", N134);
$fwrite(fileout1,"%b ", N134);
$fwrite(fileout,"N135 = %b\n", N135);
$fwrite(fileout1,"%b ", N135);
$fwrite(fileout,"N136 = %b\n", N136);
$fwrite(fileout1,"%b ", N136);
$fwrite(fileout,"N137 = %b\n", N137);
$fwrite(fileout1,"%b ", N137);
$fwrite(fileout,"N724 = %b\n", N724);
$fwrite(fileout1,"%b ", N724);
$fwrite(fileout,"N725 = %b\n", N725);
$fwrite(fileout1,"%b ", N725);
$fwrite(fileout,"N726 = %b\n", N726);
$fwrite(fileout1,"%b ", N726);
$fwrite(fileout,"N727 = %b\n", N727);
$fwrite(fileout1,"%b ", N727);
$fwrite(fileout,"N728 = %b\n", N728);
$fwrite(fileout1,"%b ", N728);
$fwrite(fileout,"N729 = %b\n", N729);
$fwrite(fileout1,"%b ", N729);
$fwrite(fileout,"N730 = %b\n", N730);
$fwrite(fileout1,"%b ", N730);
$fwrite(fileout,"N731 = %b\n", N731);
$fwrite(fileout1,"%b ", N731);
$fwrite(fileout,"N732 = %b\n", N732);
$fwrite(fileout1,"%b ", N732);
$fwrite(fileout,"N733 = %b\n", N733);
$fwrite(fileout1,"%b ", N733);
$fwrite(fileout,"N734 = %b\n", N734);
$fwrite(fileout1,"%b ", N734);
$fwrite(fileout,"N735 = %b\n", N735);
$fwrite(fileout1,"%b ", N735);
$fwrite(fileout,"N736 = %b\n", N736);
$fwrite(fileout1,"%b ", N736);
$fwrite(fileout,"N737 = %b\n", N737);
$fwrite(fileout1,"%b ", N737);
$fwrite(fileout,"N738 = %b\n", N738);
$fwrite(fileout1,"%b ", N738);
$fwrite(fileout,"N739 = %b\n", N739);
$fwrite(fileout1,"%b ", N739);
$fwrite(fileout,"N740 = %b\n", N740);
$fwrite(fileout1,"%b ", N740);
$fwrite(fileout,"N741 = %b\n", N741);
$fwrite(fileout1,"%b ", N741);
$fwrite(fileout,"N742 = %b\n", N742);
$fwrite(fileout1,"%b ", N742);
$fwrite(fileout,"N743 = %b\n", N743);
$fwrite(fileout1,"%b ", N743);
$fwrite(fileout,"N744 = %b\n", N744);
$fwrite(fileout1,"%b ", N744);
$fwrite(fileout,"N745 = %b\n", N745);
$fwrite(fileout1,"%b ", N745);
$fwrite(fileout,"N746 = %b\n", N746);
$fwrite(fileout1,"%b ", N746);
$fwrite(fileout,"N747 = %b\n", N747);
$fwrite(fileout1,"%b ", N747);
$fwrite(fileout,"N748 = %b\n", N748);
$fwrite(fileout1,"%b ", N748);
$fwrite(fileout,"N749 = %b\n", N749);
$fwrite(fileout1,"%b ", N749);
$fwrite(fileout,"N750 = %b\n", N750);
$fwrite(fileout1,"%b ", N750);
$fwrite(fileout,"N751 = %b\n", N751);
$fwrite(fileout1,"%b ", N751);
$fwrite(fileout,"N752 = %b\n", N752);
$fwrite(fileout1,"%b ", N752);
$fwrite(fileout,"N753 = %b\n", N753);
$fwrite(fileout1,"%b ", N753);
$fwrite(fileout,"N754 = %b\n", N754);
$fwrite(fileout1,"%b ", N754);
$fwrite(fileout,"N755 = %b\n", N755);
$fwrite(fileout1,"%b ", N755);
$fwrite(fileout,"Q_N724 = %b\n", Q_N724);
$fwrite(fileout1,"%b ", Q_N724);
$fwrite(fileout,"Q_N725 = %b\n", Q_N725);
$fwrite(fileout1,"%b ", Q_N725);
$fwrite(fileout,"Q_N726 = %b\n", Q_N726);
$fwrite(fileout1,"%b ", Q_N726);
$fwrite(fileout,"Q_N727 = %b\n", Q_N727);
$fwrite(fileout1,"%b ", Q_N727);
$fwrite(fileout,"Q_N728 = %b\n", Q_N728);
$fwrite(fileout1,"%b ", Q_N728);
$fwrite(fileout,"Q_N729 = %b\n", Q_N729);
$fwrite(fileout1,"%b ", Q_N729);
$fwrite(fileout,"Q_N730 = %b\n", Q_N730);
$fwrite(fileout1,"%b ", Q_N730);
$fwrite(fileout,"Q_N731 = %b\n", Q_N731);
$fwrite(fileout1,"%b ", Q_N731);
$fwrite(fileout,"Q_N732 = %b\n", Q_N732);
$fwrite(fileout1,"%b ", Q_N732);
$fwrite(fileout,"Q_N733 = %b\n", Q_N733);
$fwrite(fileout1,"%b ", Q_N733);
$fwrite(fileout,"Q_N734 = %b\n", Q_N734);
$fwrite(fileout1,"%b ", Q_N734);
$fwrite(fileout,"Q_N735 = %b\n", Q_N735);
$fwrite(fileout1,"%b ", Q_N735);
$fwrite(fileout,"Q_N736 = %b\n", Q_N736);
$fwrite(fileout1,"%b ", Q_N736);
$fwrite(fileout,"Q_N737 = %b\n", Q_N737);
$fwrite(fileout1,"%b ", Q_N737);
$fwrite(fileout,"Q_N738 = %b\n", Q_N738);
$fwrite(fileout1,"%b ", Q_N738);
$fwrite(fileout,"Q_N739 = %b\n", Q_N739);
$fwrite(fileout1,"%b ", Q_N739);
$fwrite(fileout,"Q_N740 = %b\n", Q_N740);
$fwrite(fileout1,"%b ", Q_N740);
$fwrite(fileout,"Q_N741 = %b\n", Q_N741);
$fwrite(fileout1,"%b ", Q_N741);
$fwrite(fileout,"Q_N742 = %b\n", Q_N742);
$fwrite(fileout1,"%b ", Q_N742);
$fwrite(fileout,"Q_N743 = %b\n", Q_N743);
$fwrite(fileout1,"%b ", Q_N743);
$fwrite(fileout,"Q_N744 = %b\n", Q_N744);
$fwrite(fileout1,"%b ", Q_N744);
$fwrite(fileout,"Q_N745 = %b\n", Q_N745);
$fwrite(fileout1,"%b ", Q_N745);
$fwrite(fileout,"Q_N746 = %b\n", Q_N746);
$fwrite(fileout1,"%b ", Q_N746);
$fwrite(fileout,"Q_N747 = %b\n", Q_N747);
$fwrite(fileout1,"%b ", Q_N747);
$fwrite(fileout,"Q_N748 = %b\n", Q_N748);
$fwrite(fileout1,"%b ", Q_N748);
$fwrite(fileout,"Q_N749 = %b\n", Q_N749);
$fwrite(fileout1,"%b ", Q_N749);
$fwrite(fileout,"Q_N750 = %b\n", Q_N750);
$fwrite(fileout1,"%b ", Q_N750);
$fwrite(fileout,"Q_N751 = %b\n", Q_N751);
$fwrite(fileout1,"%b ", Q_N751);
$fwrite(fileout,"Q_N752 = %b\n", Q_N752);
$fwrite(fileout1,"%b ", Q_N752);
$fwrite(fileout,"Q_N753 = %b\n", Q_N753);
$fwrite(fileout1,"%b ", Q_N753);
$fwrite(fileout,"Q_N754 = %b\n", Q_N754);
$fwrite(fileout1,"%b ", Q_N754);
$fwrite(fileout,"Q_N755 = %b\n", Q_N755);
$fwrite(fileout1,"%b ", Q_N755);
end
endmodule

