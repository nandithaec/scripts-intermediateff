library verilog;
use verilog.vl_types.all;
entity INVX4 is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end INVX4;
