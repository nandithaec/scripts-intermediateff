library verilog;
use verilog.vl_types.all;
entity BUFX2 is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end BUFX2;
