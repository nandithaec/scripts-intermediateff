library verilog;
use verilog.vl_types.all;
entity c499 is
    port(
        N1              : in     vl_logic;
        N5              : in     vl_logic;
        N9              : in     vl_logic;
        N13             : in     vl_logic;
        N17             : in     vl_logic;
        N21             : in     vl_logic;
        N25             : in     vl_logic;
        N29             : in     vl_logic;
        N33             : in     vl_logic;
        N37             : in     vl_logic;
        N41             : in     vl_logic;
        N45             : in     vl_logic;
        N49             : in     vl_logic;
        N53             : in     vl_logic;
        N57             : in     vl_logic;
        N61             : in     vl_logic;
        N65             : in     vl_logic;
        N69             : in     vl_logic;
        N73             : in     vl_logic;
        N77             : in     vl_logic;
        N81             : in     vl_logic;
        N85             : in     vl_logic;
        N89             : in     vl_logic;
        N93             : in     vl_logic;
        N97             : in     vl_logic;
        N101            : in     vl_logic;
        N105            : in     vl_logic;
        N109            : in     vl_logic;
        N113            : in     vl_logic;
        N117            : in     vl_logic;
        N121            : in     vl_logic;
        N125            : in     vl_logic;
        N129            : in     vl_logic;
        N130            : in     vl_logic;
        N131            : in     vl_logic;
        N132            : in     vl_logic;
        N133            : in     vl_logic;
        N134            : in     vl_logic;
        N135            : in     vl_logic;
        N136            : in     vl_logic;
        N137            : in     vl_logic;
        N724            : out    vl_logic;
        N725            : out    vl_logic;
        N726            : out    vl_logic;
        N727            : out    vl_logic;
        N728            : out    vl_logic;
        N729            : out    vl_logic;
        N730            : out    vl_logic;
        N731            : out    vl_logic;
        N732            : out    vl_logic;
        N733            : out    vl_logic;
        N734            : out    vl_logic;
        N735            : out    vl_logic;
        N736            : out    vl_logic;
        N737            : out    vl_logic;
        N738            : out    vl_logic;
        N739            : out    vl_logic;
        N740            : out    vl_logic;
        N741            : out    vl_logic;
        N742            : out    vl_logic;
        N743            : out    vl_logic;
        N744            : out    vl_logic;
        N745            : out    vl_logic;
        N746            : out    vl_logic;
        N747            : out    vl_logic;
        N748            : out    vl_logic;
        N749            : out    vl_logic;
        N750            : out    vl_logic;
        N751            : out    vl_logic;
        N752            : out    vl_logic;
        N753            : out    vl_logic;
        N754            : out    vl_logic;
        N755            : out    vl_logic
    );
end c499;
