
module c499 ( N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, 
        N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, 
        N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, 
        N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, 
        N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, 
        N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
  input N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57,
         N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109,
         N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135,
         N136, N137;
  output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734,
         N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745,
         N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153;

  INVX2 U1 ( .A(n46), .Y(n1) );
  INVX2 U2 ( .A(n28), .Y(n2) );
  INVX2 U3 ( .A(n39), .Y(n3) );
  INVX2 U4 ( .A(n64), .Y(n4) );
  INVX2 U5 ( .A(n35), .Y(n5) );
  INVX2 U6 ( .A(n45), .Y(n6) );
  INVX2 U7 ( .A(n30), .Y(n7) );
  INVX2 U8 ( .A(n62), .Y(n8) );
  INVX2 U9 ( .A(n70), .Y(n9) );
  INVX2 U10 ( .A(n67), .Y(n10) );
  INVX2 U11 ( .A(n32), .Y(n11) );
  INVX2 U12 ( .A(n37), .Y(n12) );
  INVX2 U13 ( .A(N49), .Y(n13) );
  INVX2 U14 ( .A(N65), .Y(n14) );
  INVX2 U15 ( .A(N117), .Y(n15) );
  XNOR2X1 U16 ( .A(N125), .B(n16), .Y(N755) );
  NAND2X1 U17 ( .A(n17), .B(n11), .Y(n16) );
  XNOR2X1 U18 ( .A(N121), .B(n18), .Y(N754) );
  NAND2X1 U19 ( .A(n17), .B(n5), .Y(n18) );
  XOR2X1 U20 ( .A(n15), .B(n19), .Y(N753) );
  NAND2X1 U21 ( .A(n17), .B(n12), .Y(n19) );
  XNOR2X1 U22 ( .A(N113), .B(n20), .Y(N752) );
  NAND2X1 U23 ( .A(n17), .B(n3), .Y(n20) );
  AND2X1 U24 ( .A(n2), .B(n21), .Y(n17) );
  XNOR2X1 U25 ( .A(N109), .B(n22), .Y(N751) );
  NAND2X1 U26 ( .A(n23), .B(n11), .Y(n22) );
  XNOR2X1 U27 ( .A(N105), .B(n24), .Y(N750) );
  NAND2X1 U28 ( .A(n23), .B(n5), .Y(n24) );
  XNOR2X1 U29 ( .A(N101), .B(n25), .Y(N749) );
  NAND2X1 U30 ( .A(n23), .B(n12), .Y(n25) );
  XNOR2X1 U31 ( .A(N97), .B(n26), .Y(N748) );
  NAND2X1 U32 ( .A(n23), .B(n3), .Y(n26) );
  AND2X1 U33 ( .A(n27), .B(n2), .Y(n23) );
  NAND3X1 U34 ( .A(n8), .B(n29), .C(n30), .Y(n28) );
  XOR2X1 U35 ( .A(N93), .B(n31), .Y(N747) );
  NOR2X1 U36 ( .A(n32), .B(n33), .Y(n31) );
  XOR2X1 U37 ( .A(N89), .B(n34), .Y(N746) );
  NOR2X1 U38 ( .A(n35), .B(n33), .Y(n34) );
  XOR2X1 U39 ( .A(N85), .B(n36), .Y(N745) );
  NOR2X1 U40 ( .A(n37), .B(n33), .Y(n36) );
  XOR2X1 U41 ( .A(N81), .B(n38), .Y(N744) );
  NOR2X1 U42 ( .A(n39), .B(n33), .Y(n38) );
  NAND3X1 U43 ( .A(n21), .B(n29), .C(n6), .Y(n33) );
  XOR2X1 U44 ( .A(N77), .B(n40), .Y(N743) );
  NOR2X1 U45 ( .A(n32), .B(n41), .Y(n40) );
  XOR2X1 U46 ( .A(N73), .B(n42), .Y(N742) );
  NOR2X1 U47 ( .A(n35), .B(n41), .Y(n42) );
  XOR2X1 U48 ( .A(N69), .B(n43), .Y(N741) );
  NOR2X1 U49 ( .A(n37), .B(n41), .Y(n43) );
  XOR2X1 U50 ( .A(N65), .B(n44), .Y(N740) );
  NOR2X1 U51 ( .A(n39), .B(n41), .Y(n44) );
  NAND3X1 U52 ( .A(n27), .B(n29), .C(n6), .Y(n41) );
  OAI21X1 U53 ( .A(n46), .B(n47), .C(n48), .Y(n29) );
  NAND2X1 U54 ( .A(n39), .B(n49), .Y(n48) );
  OAI21X1 U55 ( .A(n11), .B(n5), .C(n50), .Y(n49) );
  OAI21X1 U56 ( .A(n51), .B(n52), .C(n37), .Y(n50) );
  NAND2X1 U57 ( .A(n35), .B(n32), .Y(n47) );
  XNOR2X1 U58 ( .A(N61), .B(n53), .Y(N739) );
  NAND2X1 U59 ( .A(n54), .B(n10), .Y(n53) );
  XNOR2X1 U60 ( .A(N57), .B(n55), .Y(N738) );
  NAND2X1 U61 ( .A(n54), .B(n9), .Y(n55) );
  XNOR2X1 U62 ( .A(N53), .B(n56), .Y(N737) );
  NAND2X1 U63 ( .A(n54), .B(n8), .Y(n56) );
  XOR2X1 U64 ( .A(n13), .B(n57), .Y(N736) );
  NAND2X1 U65 ( .A(n54), .B(n7), .Y(n57) );
  AND2X1 U66 ( .A(n4), .B(n51), .Y(n54) );
  XNOR2X1 U67 ( .A(N45), .B(n58), .Y(N735) );
  NAND2X1 U68 ( .A(n59), .B(n10), .Y(n58) );
  XNOR2X1 U69 ( .A(N41), .B(n60), .Y(N734) );
  NAND2X1 U70 ( .A(n59), .B(n9), .Y(n60) );
  XNOR2X1 U71 ( .A(N37), .B(n61), .Y(N733) );
  NAND2X1 U72 ( .A(n59), .B(n8), .Y(n61) );
  XNOR2X1 U73 ( .A(N33), .B(n63), .Y(N732) );
  NAND2X1 U74 ( .A(n59), .B(n7), .Y(n63) );
  AND2X1 U75 ( .A(n52), .B(n4), .Y(n59) );
  NAND3X1 U76 ( .A(n12), .B(n65), .C(n39), .Y(n64) );
  XOR2X1 U77 ( .A(N29), .B(n66), .Y(N731) );
  NOR2X1 U78 ( .A(n67), .B(n68), .Y(n66) );
  XOR2X1 U79 ( .A(N25), .B(n69), .Y(N730) );
  NOR2X1 U80 ( .A(n70), .B(n68), .Y(n69) );
  XOR2X1 U81 ( .A(N21), .B(n71), .Y(N729) );
  NOR2X1 U82 ( .A(n62), .B(n68), .Y(n71) );
  XOR2X1 U83 ( .A(N17), .B(n72), .Y(N728) );
  NOR2X1 U84 ( .A(n30), .B(n68), .Y(n72) );
  NAND3X1 U85 ( .A(n1), .B(n65), .C(n51), .Y(n68) );
  NOR2X1 U86 ( .A(n5), .B(n32), .Y(n51) );
  XOR2X1 U87 ( .A(N13), .B(n73), .Y(N727) );
  NOR2X1 U88 ( .A(n67), .B(n74), .Y(n73) );
  XOR2X1 U89 ( .A(N9), .B(n75), .Y(N726) );
  NOR2X1 U90 ( .A(n70), .B(n74), .Y(n75) );
  XOR2X1 U91 ( .A(N5), .B(n76), .Y(N725) );
  NOR2X1 U92 ( .A(n62), .B(n74), .Y(n76) );
  XOR2X1 U93 ( .A(N1), .B(n77), .Y(N724) );
  NOR2X1 U94 ( .A(n30), .B(n74), .Y(n77) );
  NAND3X1 U95 ( .A(n1), .B(n65), .C(n52), .Y(n74) );
  NOR2X1 U96 ( .A(n11), .B(n35), .Y(n52) );
  XOR2X1 U97 ( .A(n78), .B(n79), .Y(n35) );
  XOR2X1 U98 ( .A(n80), .B(n81), .Y(n79) );
  XOR2X1 U99 ( .A(N121), .B(N105), .Y(n81) );
  XOR2X1 U100 ( .A(N89), .B(N73), .Y(n80) );
  XOR2X1 U101 ( .A(n82), .B(n83), .Y(n78) );
  XOR2X1 U102 ( .A(n84), .B(n85), .Y(n82) );
  NAND2X1 U103 ( .A(N135), .B(N137), .Y(n84) );
  XOR2X1 U104 ( .A(n86), .B(n87), .Y(n32) );
  XOR2X1 U105 ( .A(n88), .B(n89), .Y(n87) );
  XOR2X1 U106 ( .A(N125), .B(N109), .Y(n89) );
  XOR2X1 U107 ( .A(N93), .B(N77), .Y(n88) );
  XOR2X1 U108 ( .A(n90), .B(n91), .Y(n86) );
  XOR2X1 U109 ( .A(n92), .B(n93), .Y(n90) );
  NAND2X1 U110 ( .A(N136), .B(N137), .Y(n92) );
  OAI21X1 U111 ( .A(n45), .B(n94), .C(n95), .Y(n65) );
  NAND2X1 U112 ( .A(n30), .B(n96), .Y(n95) );
  OAI21X1 U113 ( .A(n9), .B(n10), .C(n97), .Y(n96) );
  OAI21X1 U114 ( .A(n21), .B(n27), .C(n62), .Y(n97) );
  NOR2X1 U115 ( .A(n10), .B(n70), .Y(n27) );
  NOR2X1 U116 ( .A(n9), .B(n67), .Y(n21) );
  NAND2X1 U117 ( .A(n70), .B(n67), .Y(n94) );
  XOR2X1 U118 ( .A(n98), .B(n99), .Y(n67) );
  XOR2X1 U119 ( .A(n100), .B(n101), .Y(n99) );
  XOR2X1 U120 ( .A(N29), .B(N13), .Y(n101) );
  XOR2X1 U121 ( .A(N61), .B(N45), .Y(n100) );
  XOR2X1 U122 ( .A(n102), .B(n103), .Y(n98) );
  XOR2X1 U123 ( .A(n104), .B(n105), .Y(n102) );
  NAND2X1 U124 ( .A(N132), .B(N137), .Y(n104) );
  XOR2X1 U125 ( .A(n106), .B(n107), .Y(n70) );
  XOR2X1 U126 ( .A(n108), .B(n109), .Y(n107) );
  XOR2X1 U127 ( .A(N41), .B(N25), .Y(n109) );
  XOR2X1 U128 ( .A(N9), .B(N57), .Y(n108) );
  XOR2X1 U129 ( .A(n110), .B(n111), .Y(n106) );
  XOR2X1 U130 ( .A(n112), .B(n113), .Y(n110) );
  NAND2X1 U131 ( .A(N131), .B(N137), .Y(n112) );
  NAND2X1 U132 ( .A(n62), .B(n7), .Y(n45) );
  XOR2X1 U133 ( .A(n114), .B(n115), .Y(n62) );
  XOR2X1 U134 ( .A(n116), .B(n117), .Y(n115) );
  XOR2X1 U135 ( .A(N37), .B(N21), .Y(n117) );
  XOR2X1 U136 ( .A(N53), .B(N5), .Y(n116) );
  XOR2X1 U137 ( .A(n118), .B(n111), .Y(n114) );
  XNOR2X1 U138 ( .A(n119), .B(n120), .Y(n111) );
  XOR2X1 U139 ( .A(N97), .B(N109), .Y(n120) );
  XNOR2X1 U140 ( .A(N101), .B(N105), .Y(n119) );
  XOR2X1 U141 ( .A(n121), .B(n103), .Y(n118) );
  XNOR2X1 U142 ( .A(n122), .B(n123), .Y(n103) );
  XOR2X1 U143 ( .A(N125), .B(N121), .Y(n123) );
  XOR2X1 U144 ( .A(N113), .B(n15), .Y(n122) );
  NAND2X1 U145 ( .A(N130), .B(N137), .Y(n121) );
  NAND2X1 U146 ( .A(n37), .B(n3), .Y(n46) );
  XOR2X1 U147 ( .A(n124), .B(n125), .Y(n39) );
  XOR2X1 U148 ( .A(n126), .B(n127), .Y(n125) );
  XOR2X1 U149 ( .A(N65), .B(N113), .Y(n127) );
  XOR2X1 U150 ( .A(N97), .B(N81), .Y(n126) );
  XOR2X1 U151 ( .A(n128), .B(n85), .Y(n124) );
  XNOR2X1 U152 ( .A(n129), .B(n130), .Y(n85) );
  XOR2X1 U153 ( .A(N9), .B(N5), .Y(n130) );
  XNOR2X1 U154 ( .A(N1), .B(N13), .Y(n129) );
  XOR2X1 U155 ( .A(n131), .B(n93), .Y(n128) );
  XNOR2X1 U156 ( .A(n132), .B(n133), .Y(n93) );
  XOR2X1 U157 ( .A(N29), .B(N25), .Y(n133) );
  XNOR2X1 U158 ( .A(N17), .B(N21), .Y(n132) );
  NAND2X1 U159 ( .A(N133), .B(N137), .Y(n131) );
  XOR2X1 U160 ( .A(n134), .B(n135), .Y(n37) );
  XOR2X1 U161 ( .A(n136), .B(n137), .Y(n135) );
  XOR2X1 U162 ( .A(N117), .B(N101), .Y(n137) );
  XOR2X1 U163 ( .A(N85), .B(N69), .Y(n136) );
  XOR2X1 U164 ( .A(n138), .B(n83), .Y(n134) );
  XNOR2X1 U165 ( .A(n139), .B(n140), .Y(n83) );
  XOR2X1 U166 ( .A(N45), .B(N41), .Y(n140) );
  XNOR2X1 U167 ( .A(N33), .B(N37), .Y(n139) );
  XOR2X1 U168 ( .A(n141), .B(n91), .Y(n138) );
  XNOR2X1 U169 ( .A(n142), .B(n143), .Y(n91) );
  XOR2X1 U170 ( .A(N61), .B(N57), .Y(n143) );
  XOR2X1 U171 ( .A(n13), .B(N53), .Y(n142) );
  NAND2X1 U172 ( .A(N137), .B(N134), .Y(n141) );
  XOR2X1 U173 ( .A(n144), .B(n145), .Y(n30) );
  XOR2X1 U174 ( .A(n146), .B(n147), .Y(n145) );
  XOR2X1 U175 ( .A(N17), .B(N1), .Y(n147) );
  XOR2X1 U176 ( .A(N49), .B(N33), .Y(n146) );
  XOR2X1 U177 ( .A(n148), .B(n113), .Y(n144) );
  XNOR2X1 U178 ( .A(n149), .B(n150), .Y(n113) );
  XOR2X1 U179 ( .A(N77), .B(N73), .Y(n150) );
  XOR2X1 U180 ( .A(n14), .B(N69), .Y(n149) );
  XOR2X1 U181 ( .A(n151), .B(n105), .Y(n148) );
  XNOR2X1 U182 ( .A(n152), .B(n153), .Y(n105) );
  XOR2X1 U183 ( .A(N93), .B(N89), .Y(n153) );
  XNOR2X1 U184 ( .A(N81), .B(N85), .Y(n152) );
  NAND2X1 U185 ( .A(N129), .B(N137), .Y(n151) );
endmodule


module dff_104 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_103 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_102 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_101 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_100 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_99 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_98 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_97 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_96 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_95 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_94 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_93 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_92 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_91 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_90 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_89 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_88 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_87 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_86 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_85 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_84 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_83 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_82 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_81 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_80 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_79 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_78 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_77 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_76 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_75 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_74 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_73 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_72 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_71 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_70 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_69 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_68 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_67 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_66 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_65 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_64 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_63 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_62 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_61 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_60 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_59 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_58 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_57 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_56 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_55 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_54 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_53 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_52 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_51 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_50 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_49 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_48 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_47 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_46 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_45 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_44 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_43 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_42 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_41 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_40 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_39 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_38 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_37 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_36 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_35 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_34 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_33 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_32 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_31 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_30 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_29 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_28 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_27 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_26 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_25 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_24 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_23 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_22 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_21 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_20 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_19 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_18 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_17 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_16 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_15 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_14 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_13 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_12 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_11 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_10 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_9 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_8 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_7 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_6 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_5 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_4 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_3 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_2 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_1 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_0 ( q, d, clk );
  input d, clk;
  output q;


  DFFPOSX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module c499_clk_opFF ( clk, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, 
        N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, 
        N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, 
        N134, N135, N136, N137, Qout_N724, Qout_N725, Qout_N726, Qout_N727, 
        Qout_N728, Qout_N729, Qout_N730, Qout_N731, Qout_N732, Qout_N733, 
        Qout_N734, Qout_N735, Qout_N736, Qout_N737, Qout_N738, Qout_N739, 
        Qout_N740, Qout_N741, Qout_N742, Qout_N743, Qout_N744, Qout_N745, 
        Qout_N746, Qout_N747, Qout_N748, Qout_N749, Qout_N750, Qout_N751, 
        Qout_N752, Qout_N753, Qout_N754, Qout_N755 );
  input clk, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53,
         N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105,
         N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134,
         N135, N136, N137;
  output Qout_N724, Qout_N725, Qout_N726, Qout_N727, Qout_N728, Qout_N729,
         Qout_N730, Qout_N731, Qout_N732, Qout_N733, Qout_N734, Qout_N735,
         Qout_N736, Qout_N737, Qout_N738, Qout_N739, Qout_N740, Qout_N741,
         Qout_N742, Qout_N743, Qout_N744, Qout_N745, Qout_N746, Qout_N747,
         Qout_N748, Qout_N749, Qout_N750, Qout_N751, Qout_N752, Qout_N753,
         Qout_N754, Qout_N755;
  wire   IN_N1, IN_N5, IN_N9, IN_N13, IN_N17, IN_N21, IN_N25, IN_N29, IN_N33,
         IN_N37, IN_N41, IN_N45, IN_N49, IN_N53, IN_N57, IN_N61, IN_N65,
         IN_N69, IN_N73, IN_N77, IN_N81, IN_N85, IN_N89, IN_N93, IN_N97,
         IN_N101, IN_N105, IN_N109, IN_N113, IN_N117, IN_N121, IN_N125,
         IN_N129, IN_N130, IN_N131, IN_N132, IN_N133, IN_N134, IN_N135,
         IN_N136, IN_N137, N724, N725, N726, N727, N728, N729, N730, N731,
         N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742,
         N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753,
         N754, N755, Q_N724, Q_N725, Q_N726, Q_N727, Q_N728, Q_N729, Q_N730,
         Q_N731, Q_N732, Q_N733, Q_N734, Q_N735, Q_N736, Q_N737, Q_N738,
         Q_N739, Q_N740, Q_N741, Q_N742, Q_N743, Q_N744, Q_N745, Q_N746,
         Q_N747, Q_N748, Q_N749, Q_N750, Q_N751, Q_N752, Q_N753, Q_N754,
         Q_N755;

  c499 c0 ( .N1(IN_N1), .N5(IN_N5), .N9(IN_N9), .N13(IN_N13), .N17(IN_N17), 
        .N21(IN_N21), .N25(IN_N25), .N29(IN_N29), .N33(IN_N33), .N37(IN_N37), 
        .N41(IN_N41), .N45(IN_N45), .N49(IN_N49), .N53(IN_N53), .N57(IN_N57), 
        .N61(IN_N61), .N65(IN_N65), .N69(IN_N69), .N73(IN_N73), .N77(IN_N77), 
        .N81(IN_N81), .N85(IN_N85), .N89(IN_N89), .N93(IN_N93), .N97(IN_N97), 
        .N101(IN_N101), .N105(IN_N105), .N109(IN_N109), .N113(IN_N113), .N117(
        IN_N117), .N121(IN_N121), .N125(IN_N125), .N129(IN_N129), .N130(
        IN_N130), .N131(IN_N131), .N132(IN_N132), .N133(IN_N133), .N134(
        IN_N134), .N135(IN_N135), .N136(IN_N136), .N137(IN_N137), .N724(N724), 
        .N725(N725), .N726(N726), .N727(N727), .N728(N728), .N729(N729), 
        .N730(N730), .N731(N731), .N732(N732), .N733(N733), .N734(N734), 
        .N735(N735), .N736(N736), .N737(N737), .N738(N738), .N739(N739), 
        .N740(N740), .N741(N741), .N742(N742), .N743(N743), .N744(N744), 
        .N745(N745), .N746(N746), .N747(N747), .N748(N748), .N749(N749), 
        .N750(N750), .N751(N751), .N752(N752), .N753(N753), .N754(N754), 
        .N755(N755) );
  dff_104 iDFF_1 ( .q(IN_N1), .d(N1), .clk(clk) );
  dff_103 iDFF_2 ( .q(IN_N5), .d(N5), .clk(clk) );
  dff_102 iDFF_3 ( .q(IN_N9), .d(N9), .clk(clk) );
  dff_101 iDFF_4 ( .q(IN_N13), .d(N13), .clk(clk) );
  dff_100 iDFF_5 ( .q(IN_N17), .d(N17), .clk(clk) );
  dff_99 iDFF_6 ( .q(IN_N21), .d(N21), .clk(clk) );
  dff_98 iDFF_7 ( .q(IN_N25), .d(N25), .clk(clk) );
  dff_97 iDFF_8 ( .q(IN_N29), .d(N29), .clk(clk) );
  dff_96 iDFF_9 ( .q(IN_N33), .d(N33), .clk(clk) );
  dff_95 iDFF_10 ( .q(IN_N37), .d(N37), .clk(clk) );
  dff_94 iDFF_11 ( .q(IN_N41), .d(N41), .clk(clk) );
  dff_93 iDFF_12 ( .q(IN_N45), .d(N45), .clk(clk) );
  dff_92 iDFF_13 ( .q(IN_N49), .d(N49), .clk(clk) );
  dff_91 iDFF_14 ( .q(IN_N53), .d(N53), .clk(clk) );
  dff_90 iDFF_15 ( .q(IN_N57), .d(N57), .clk(clk) );
  dff_89 iDFF_16 ( .q(IN_N61), .d(N61), .clk(clk) );
  dff_88 iDFF_17 ( .q(IN_N65), .d(N65), .clk(clk) );
  dff_87 iDFF_18 ( .q(IN_N69), .d(N69), .clk(clk) );
  dff_86 iDFF_19 ( .q(IN_N73), .d(N73), .clk(clk) );
  dff_85 iDFF_20 ( .q(IN_N77), .d(N77), .clk(clk) );
  dff_84 iDFF_21 ( .q(IN_N81), .d(N81), .clk(clk) );
  dff_83 iDFF_22 ( .q(IN_N85), .d(N85), .clk(clk) );
  dff_82 iDFF_23 ( .q(IN_N89), .d(N89), .clk(clk) );
  dff_81 iDFF_24 ( .q(IN_N93), .d(N93), .clk(clk) );
  dff_80 iDFF_25 ( .q(IN_N97), .d(N97), .clk(clk) );
  dff_79 iDFF_26 ( .q(IN_N101), .d(N101), .clk(clk) );
  dff_78 iDFF_27 ( .q(IN_N105), .d(N105), .clk(clk) );
  dff_77 iDFF_28 ( .q(IN_N109), .d(N109), .clk(clk) );
  dff_76 iDFF_29 ( .q(IN_N113), .d(N113), .clk(clk) );
  dff_75 iDFF_30 ( .q(IN_N117), .d(N117), .clk(clk) );
  dff_74 iDFF_31 ( .q(IN_N121), .d(N121), .clk(clk) );
  dff_73 iDFF_32 ( .q(IN_N125), .d(N125), .clk(clk) );
  dff_72 iDFF_33 ( .q(IN_N129), .d(N129), .clk(clk) );
  dff_71 iDFF_34 ( .q(IN_N130), .d(N130), .clk(clk) );
  dff_70 iDFF_35 ( .q(IN_N131), .d(N131), .clk(clk) );
  dff_69 iDFF_36 ( .q(IN_N132), .d(N132), .clk(clk) );
  dff_68 iDFF_37 ( .q(IN_N133), .d(N133), .clk(clk) );
  dff_67 iDFF_38 ( .q(IN_N134), .d(N134), .clk(clk) );
  dff_66 iDFF_39 ( .q(IN_N135), .d(N135), .clk(clk) );
  dff_65 iDFF_40 ( .q(IN_N136), .d(N136), .clk(clk) );
  dff_64 iDFF_41 ( .q(IN_N137), .d(N137), .clk(clk) );
  dff_63 DFF_1 ( .q(Q_N724), .d(N724), .clk(clk) );
  dff_62 DFF_2 ( .q(Q_N725), .d(N725), .clk(clk) );
  dff_61 DFF_3 ( .q(Q_N726), .d(N726), .clk(clk) );
  dff_60 DFF_4 ( .q(Q_N727), .d(N727), .clk(clk) );
  dff_59 DFF_5 ( .q(Q_N728), .d(N728), .clk(clk) );
  dff_58 DFF_6 ( .q(Q_N729), .d(N729), .clk(clk) );
  dff_57 DFF_7 ( .q(Q_N730), .d(N730), .clk(clk) );
  dff_56 DFF_8 ( .q(Q_N731), .d(N731), .clk(clk) );
  dff_55 DFF_9 ( .q(Q_N732), .d(N732), .clk(clk) );
  dff_54 DFF_10 ( .q(Q_N733), .d(N733), .clk(clk) );
  dff_53 DFF_11 ( .q(Q_N734), .d(N734), .clk(clk) );
  dff_52 DFF_12 ( .q(Q_N735), .d(N735), .clk(clk) );
  dff_51 DFF_13 ( .q(Q_N736), .d(N736), .clk(clk) );
  dff_50 DFF_14 ( .q(Q_N737), .d(N737), .clk(clk) );
  dff_49 DFF_15 ( .q(Q_N738), .d(N738), .clk(clk) );
  dff_48 DFF_16 ( .q(Q_N739), .d(N739), .clk(clk) );
  dff_47 DFF_17 ( .q(Q_N740), .d(N740), .clk(clk) );
  dff_46 DFF_18 ( .q(Q_N741), .d(N741), .clk(clk) );
  dff_45 DFF_19 ( .q(Q_N742), .d(N742), .clk(clk) );
  dff_44 DFF_20 ( .q(Q_N743), .d(N743), .clk(clk) );
  dff_43 DFF_21 ( .q(Q_N744), .d(N744), .clk(clk) );
  dff_42 DFF_22 ( .q(Q_N745), .d(N745), .clk(clk) );
  dff_41 DFF_23 ( .q(Q_N746), .d(N746), .clk(clk) );
  dff_40 DFF_24 ( .q(Q_N747), .d(N747), .clk(clk) );
  dff_39 DFF_25 ( .q(Q_N748), .d(N748), .clk(clk) );
  dff_38 DFF_26 ( .q(Q_N749), .d(N749), .clk(clk) );
  dff_37 DFF_27 ( .q(Q_N750), .d(N750), .clk(clk) );
  dff_36 DFF_28 ( .q(Q_N751), .d(N751), .clk(clk) );
  dff_35 DFF_29 ( .q(Q_N752), .d(N752), .clk(clk) );
  dff_34 DFF_30 ( .q(Q_N753), .d(N753), .clk(clk) );
  dff_33 DFF_31 ( .q(Q_N754), .d(N754), .clk(clk) );
  dff_32 DFF_32 ( .q(Q_N755), .d(N755), .clk(clk) );
  dff_31 oDFF_1 ( .q(Qout_N724), .d(Q_N724), .clk(clk) );
  dff_30 oDFF_2 ( .q(Qout_N725), .d(Q_N725), .clk(clk) );
  dff_29 oDFF_3 ( .q(Qout_N726), .d(Q_N726), .clk(clk) );
  dff_28 oDFF_4 ( .q(Qout_N727), .d(Q_N727), .clk(clk) );
  dff_27 oDFF_5 ( .q(Qout_N728), .d(Q_N728), .clk(clk) );
  dff_26 oDFF_6 ( .q(Qout_N729), .d(Q_N729), .clk(clk) );
  dff_25 oDFF_7 ( .q(Qout_N730), .d(Q_N730), .clk(clk) );
  dff_24 oDFF_8 ( .q(Qout_N731), .d(Q_N731), .clk(clk) );
  dff_23 oDFF_9 ( .q(Qout_N732), .d(Q_N732), .clk(clk) );
  dff_22 oDFF_10 ( .q(Qout_N733), .d(Q_N733), .clk(clk) );
  dff_21 oDFF_11 ( .q(Qout_N734), .d(Q_N734), .clk(clk) );
  dff_20 oDFF_12 ( .q(Qout_N735), .d(Q_N735), .clk(clk) );
  dff_19 oDFF_13 ( .q(Qout_N736), .d(Q_N736), .clk(clk) );
  dff_18 oDFF_14 ( .q(Qout_N737), .d(Q_N737), .clk(clk) );
  dff_17 oDFF_15 ( .q(Qout_N738), .d(Q_N738), .clk(clk) );
  dff_16 oDFF_16 ( .q(Qout_N739), .d(Q_N739), .clk(clk) );
  dff_15 oDFF_17 ( .q(Qout_N740), .d(Q_N740), .clk(clk) );
  dff_14 oDFF_18 ( .q(Qout_N741), .d(Q_N741), .clk(clk) );
  dff_13 oDFF_19 ( .q(Qout_N742), .d(Q_N742), .clk(clk) );
  dff_12 oDFF_20 ( .q(Qout_N743), .d(Q_N743), .clk(clk) );
  dff_11 oDFF_21 ( .q(Qout_N744), .d(Q_N744), .clk(clk) );
  dff_10 oDFF_22 ( .q(Qout_N745), .d(Q_N745), .clk(clk) );
  dff_9 oDFF_23 ( .q(Qout_N746), .d(Q_N746), .clk(clk) );
  dff_8 oDFF_24 ( .q(Qout_N747), .d(Q_N747), .clk(clk) );
  dff_7 oDFF_25 ( .q(Qout_N748), .d(Q_N748), .clk(clk) );
  dff_6 oDFF_26 ( .q(Qout_N749), .d(Q_N749), .clk(clk) );
  dff_5 oDFF_27 ( .q(Qout_N750), .d(Q_N750), .clk(clk) );
  dff_4 oDFF_28 ( .q(Qout_N751), .d(Q_N751), .clk(clk) );
  dff_3 oDFF_29 ( .q(Qout_N752), .d(Q_N752), .clk(clk) );
  dff_2 oDFF_30 ( .q(Qout_N753), .d(Q_N753), .clk(clk) );
  dff_1 oDFF_31 ( .q(Qout_N754), .d(Q_N754), .clk(clk) );
  dff_0 oDFF_32 ( .q(Qout_N755), .d(Q_N755), .clk(clk) );
endmodule

