
library IEEE;

use IEEE.std_logic_1164.all;

entity dff_103 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_103;

architecture SYN_verilog of dff_103 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_102 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_102;

architecture SYN_verilog of dff_102 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_101 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_101;

architecture SYN_verilog of dff_101 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_100 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_100;

architecture SYN_verilog of dff_100 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_99 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_99;

architecture SYN_verilog of dff_99 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_98 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_98;

architecture SYN_verilog of dff_98 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_97 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_97;

architecture SYN_verilog of dff_97 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_96 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_96;

architecture SYN_verilog of dff_96 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_95 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_95;

architecture SYN_verilog of dff_95 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_94 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_94;

architecture SYN_verilog of dff_94 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_93 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_93;

architecture SYN_verilog of dff_93 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_92 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_92;

architecture SYN_verilog of dff_92 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_91 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_91;

architecture SYN_verilog of dff_91 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_90 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_90;

architecture SYN_verilog of dff_90 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_89 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_89;

architecture SYN_verilog of dff_89 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_88 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_88;

architecture SYN_verilog of dff_88 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_87 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_87;

architecture SYN_verilog of dff_87 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_86 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_86;

architecture SYN_verilog of dff_86 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_85 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_85;

architecture SYN_verilog of dff_85 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_84 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_84;

architecture SYN_verilog of dff_84 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_83 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_83;

architecture SYN_verilog of dff_83 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_82 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_82;

architecture SYN_verilog of dff_82 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_81 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_81;

architecture SYN_verilog of dff_81 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_80 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_80;

architecture SYN_verilog of dff_80 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_79 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_79;

architecture SYN_verilog of dff_79 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_78 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_78;

architecture SYN_verilog of dff_78 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_77 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_77;

architecture SYN_verilog of dff_77 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_76 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_76;

architecture SYN_verilog of dff_76 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_75 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_75;

architecture SYN_verilog of dff_75 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_74 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_74;

architecture SYN_verilog of dff_74 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_73 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_73;

architecture SYN_verilog of dff_73 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_72 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_72;

architecture SYN_verilog of dff_72 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_71 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_71;

architecture SYN_verilog of dff_71 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_70 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_70;

architecture SYN_verilog of dff_70 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_69 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_69;

architecture SYN_verilog of dff_69 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_68 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_68;

architecture SYN_verilog of dff_68 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_67 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_67;

architecture SYN_verilog of dff_67 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_66 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_66;

architecture SYN_verilog of dff_66 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_65 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_65;

architecture SYN_verilog of dff_65 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_64 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_64;

architecture SYN_verilog of dff_64 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_63 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_63;

architecture SYN_verilog of dff_63 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_62 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_62;

architecture SYN_verilog of dff_62 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_61 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_61;

architecture SYN_verilog of dff_61 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_60 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_60;

architecture SYN_verilog of dff_60 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_59 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_59;

architecture SYN_verilog of dff_59 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_58 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_58;

architecture SYN_verilog of dff_58 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_57 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_57;

architecture SYN_verilog of dff_57 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_56 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_56;

architecture SYN_verilog of dff_56 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_55 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_55;

architecture SYN_verilog of dff_55 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_54 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_54;

architecture SYN_verilog of dff_54 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_53 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_53;

architecture SYN_verilog of dff_53 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_52 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_52;

architecture SYN_verilog of dff_52 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_51 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_51;

architecture SYN_verilog of dff_51 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_50 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_50;

architecture SYN_verilog of dff_50 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_49 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_49;

architecture SYN_verilog of dff_49 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_48 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_48;

architecture SYN_verilog of dff_48 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_47 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_47;

architecture SYN_verilog of dff_47 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_46 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_46;

architecture SYN_verilog of dff_46 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_45 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_45;

architecture SYN_verilog of dff_45 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_44 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_44;

architecture SYN_verilog of dff_44 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_43 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_43;

architecture SYN_verilog of dff_43 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_42 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_42;

architecture SYN_verilog of dff_42 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_41 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_41;

architecture SYN_verilog of dff_41 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_40 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_40;

architecture SYN_verilog of dff_40 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_39 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_39;

architecture SYN_verilog of dff_39 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_38 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_38;

architecture SYN_verilog of dff_38 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_37 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_37;

architecture SYN_verilog of dff_37 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_36 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_36;

architecture SYN_verilog of dff_36 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_35 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_35;

architecture SYN_verilog of dff_35 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_34 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_34;

architecture SYN_verilog of dff_34 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_33 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_33;

architecture SYN_verilog of dff_33 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_32 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_32;

architecture SYN_verilog of dff_32 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_31 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_31;

architecture SYN_verilog of dff_31 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_30 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_30;

architecture SYN_verilog of dff_30 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_29 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_29;

architecture SYN_verilog of dff_29 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_28 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_28;

architecture SYN_verilog of dff_28 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_27 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_27;

architecture SYN_verilog of dff_27 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_26 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_26;

architecture SYN_verilog of dff_26 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_25 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_25;

architecture SYN_verilog of dff_25 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_24 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_24;

architecture SYN_verilog of dff_24 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_23 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_23;

architecture SYN_verilog of dff_23 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_22 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_22;

architecture SYN_verilog of dff_22 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_21 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_21;

architecture SYN_verilog of dff_21 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_20 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_20;

architecture SYN_verilog of dff_20 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_19 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_19;

architecture SYN_verilog of dff_19 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_18 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_18;

architecture SYN_verilog of dff_18 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_17 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_17;

architecture SYN_verilog of dff_17 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_16 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_16;

architecture SYN_verilog of dff_16 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_15 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_15;

architecture SYN_verilog of dff_15 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_14 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_14;

architecture SYN_verilog of dff_14 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_13 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_13;

architecture SYN_verilog of dff_13 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_12 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_12;

architecture SYN_verilog of dff_12 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_11 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_11;

architecture SYN_verilog of dff_11 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_10 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_10;

architecture SYN_verilog of dff_10 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_9 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_9;

architecture SYN_verilog of dff_9 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_8 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_8;

architecture SYN_verilog of dff_8 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_7 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_7;

architecture SYN_verilog of dff_7 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_6 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_6;

architecture SYN_verilog of dff_6 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_5 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_5;

architecture SYN_verilog of dff_5 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_4 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_4;

architecture SYN_verilog of dff_4 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_3 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_3;

architecture SYN_verilog of dff_3 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_2 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_2;

architecture SYN_verilog of dff_2 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_1 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_1;

architecture SYN_verilog of dff_1 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_0 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_0;

architecture SYN_verilog of dff_0 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity dff_104 is

   port( q : out std_logic;  d, clk : in std_logic);

end dff_104;

architecture SYN_verilog of dff_104 is

   component DFFPOSX1
      port( D, CLK : in std_logic;  Q : out std_logic);
   end component;

begin
   
   q_reg : DFFPOSX1 port map( D => d, CLK => clk, Q => q);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity c499 is

   port( N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57
         , N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, 
         N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136
         , N137 : in std_logic;  N724, N725, N726, N727, N728, N729, N730, N731
         , N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, 
         N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754
         , N755 : out std_logic);

end c499;

architecture SYN_verilog of c499 is

   component NAND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XNOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component XOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component NOR2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component OAI21X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component NAND3X1
      port( A, B, C : in std_logic;  Y : out std_logic);
   end component;
   
   component AND2X1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component INVX2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1_port, n2, n3, n4, n5_port, n6, n7, n8, n9_port, n10, n11, n12, 
      n13_port, n14, n15, n16, n17_port, n18, n19, n20, n21_port, n22, n23, n24
      , n25_port, n26, n27, n28, n29_port, n30, n31, n32, n33_port, n34, n35, 
      n36, n37_port, n38, n39, n40, n41_port, n42, n43, n44, n45_port, n46, n47
      , n48, n49_port, n50, n51, n52, n53_port, n54, n55, n56, n57_port, n58, 
      n59, n60, n61_port, n62, n63, n64, n65_port, n66, n67, n68, n69_port, n70
      , n71, n72, n73_port, n74, n75, n76, n77_port, n78, n79, n80, n81_port, 
      n82, n83, n84, n85_port, n86, n87, n88, n89_port, n90, n91, n92, n93_port
      , n94, n95, n96, n97_port, n98, n99, n100, n101_port, n102, n103, n104, 
      n105_port, n106, n107, n108, n109_port, n110, n111, n112, n113_port, n114
      , n115, n116, n117_port, n118, n119, n120, n121_port, n122, n123, n124, 
      n125_port, n126, n127, n128, n129_port, n130_port, n131_port, n132_port, 
      n133_port, n134_port, n135_port, n136_port, n137_port, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153 : std_logic;

begin
   
   U1 : INVX2 port map( A => n46, Y => n1_port);
   U2 : INVX2 port map( A => n28, Y => n2);
   U3 : INVX2 port map( A => n39, Y => n3);
   U4 : INVX2 port map( A => n64, Y => n4);
   U5 : INVX2 port map( A => n35, Y => n5_port);
   U6 : INVX2 port map( A => n45_port, Y => n6);
   U7 : INVX2 port map( A => n30, Y => n7);
   U8 : INVX2 port map( A => n62, Y => n8);
   U9 : INVX2 port map( A => n70, Y => n9_port);
   U10 : INVX2 port map( A => n67, Y => n10);
   U11 : INVX2 port map( A => n32, Y => n11);
   U12 : INVX2 port map( A => n37_port, Y => n12);
   U13 : INVX2 port map( A => N49, Y => n13_port);
   U14 : INVX2 port map( A => N65, Y => n14);
   U15 : INVX2 port map( A => N117, Y => n15);
   U16 : XNOR2X1 port map( A => N125, B => n16, Y => N755);
   U17 : NAND2X1 port map( A => n17_port, B => n11, Y => n16);
   U18 : XNOR2X1 port map( A => N121, B => n18, Y => N754);
   U19 : NAND2X1 port map( A => n17_port, B => n5_port, Y => n18);
   U20 : XOR2X1 port map( A => n15, B => n19, Y => N753);
   U21 : NAND2X1 port map( A => n17_port, B => n12, Y => n19);
   U22 : XNOR2X1 port map( A => N113, B => n20, Y => N752);
   U23 : NAND2X1 port map( A => n17_port, B => n3, Y => n20);
   U24 : AND2X1 port map( A => n2, B => n21_port, Y => n17_port);
   U25 : XNOR2X1 port map( A => N109, B => n22, Y => N751);
   U26 : NAND2X1 port map( A => n23, B => n11, Y => n22);
   U27 : XNOR2X1 port map( A => N105, B => n24, Y => N750);
   U28 : NAND2X1 port map( A => n23, B => n5_port, Y => n24);
   U29 : XNOR2X1 port map( A => N101, B => n25_port, Y => N749);
   U30 : NAND2X1 port map( A => n23, B => n12, Y => n25_port);
   U31 : XNOR2X1 port map( A => N97, B => n26, Y => N748);
   U32 : NAND2X1 port map( A => n23, B => n3, Y => n26);
   U33 : AND2X1 port map( A => n27, B => n2, Y => n23);
   U34 : NAND3X1 port map( A => n8, B => n29_port, C => n30, Y => n28);
   U35 : XOR2X1 port map( A => N93, B => n31, Y => N747);
   U36 : NOR2X1 port map( A => n32, B => n33_port, Y => n31);
   U37 : XOR2X1 port map( A => N89, B => n34, Y => N746);
   U38 : NOR2X1 port map( A => n35, B => n33_port, Y => n34);
   U39 : XOR2X1 port map( A => N85, B => n36, Y => N745);
   U40 : NOR2X1 port map( A => n37_port, B => n33_port, Y => n36);
   U41 : XOR2X1 port map( A => N81, B => n38, Y => N744);
   U42 : NOR2X1 port map( A => n39, B => n33_port, Y => n38);
   U43 : NAND3X1 port map( A => n21_port, B => n29_port, C => n6, Y => n33_port
                           );
   U44 : XOR2X1 port map( A => N77, B => n40, Y => N743);
   U45 : NOR2X1 port map( A => n32, B => n41_port, Y => n40);
   U46 : XOR2X1 port map( A => N73, B => n42, Y => N742);
   U47 : NOR2X1 port map( A => n35, B => n41_port, Y => n42);
   U48 : XOR2X1 port map( A => N69, B => n43, Y => N741);
   U49 : NOR2X1 port map( A => n37_port, B => n41_port, Y => n43);
   U50 : XOR2X1 port map( A => N65, B => n44, Y => N740);
   U51 : NOR2X1 port map( A => n39, B => n41_port, Y => n44);
   U52 : NAND3X1 port map( A => n27, B => n29_port, C => n6, Y => n41_port);
   U53 : OAI21X1 port map( A => n46, B => n47, C => n48, Y => n29_port);
   U54 : NAND2X1 port map( A => n39, B => n49_port, Y => n48);
   U55 : OAI21X1 port map( A => n11, B => n5_port, C => n50, Y => n49_port);
   U56 : OAI21X1 port map( A => n51, B => n52, C => n37_port, Y => n50);
   U57 : NAND2X1 port map( A => n35, B => n32, Y => n47);
   U58 : XNOR2X1 port map( A => N61, B => n53_port, Y => N739);
   U59 : NAND2X1 port map( A => n54, B => n10, Y => n53_port);
   U60 : XNOR2X1 port map( A => N57, B => n55, Y => N738);
   U61 : NAND2X1 port map( A => n54, B => n9_port, Y => n55);
   U62 : XNOR2X1 port map( A => N53, B => n56, Y => N737);
   U63 : NAND2X1 port map( A => n54, B => n8, Y => n56);
   U64 : XOR2X1 port map( A => n13_port, B => n57_port, Y => N736);
   U65 : NAND2X1 port map( A => n54, B => n7, Y => n57_port);
   U66 : AND2X1 port map( A => n4, B => n51, Y => n54);
   U67 : XNOR2X1 port map( A => N45, B => n58, Y => N735);
   U68 : NAND2X1 port map( A => n59, B => n10, Y => n58);
   U69 : XNOR2X1 port map( A => N41, B => n60, Y => N734);
   U70 : NAND2X1 port map( A => n59, B => n9_port, Y => n60);
   U71 : XNOR2X1 port map( A => N37, B => n61_port, Y => N733);
   U72 : NAND2X1 port map( A => n59, B => n8, Y => n61_port);
   U73 : XNOR2X1 port map( A => N33, B => n63, Y => N732);
   U74 : NAND2X1 port map( A => n59, B => n7, Y => n63);
   U75 : AND2X1 port map( A => n52, B => n4, Y => n59);
   U76 : NAND3X1 port map( A => n12, B => n65_port, C => n39, Y => n64);
   U77 : XOR2X1 port map( A => N29, B => n66, Y => N731);
   U78 : NOR2X1 port map( A => n67, B => n68, Y => n66);
   U79 : XOR2X1 port map( A => N25, B => n69_port, Y => N730);
   U80 : NOR2X1 port map( A => n70, B => n68, Y => n69_port);
   U81 : XOR2X1 port map( A => N21, B => n71, Y => N729);
   U82 : NOR2X1 port map( A => n62, B => n68, Y => n71);
   U83 : XOR2X1 port map( A => N17, B => n72, Y => N728);
   U84 : NOR2X1 port map( A => n30, B => n68, Y => n72);
   U85 : NAND3X1 port map( A => n1_port, B => n65_port, C => n51, Y => n68);
   U86 : NOR2X1 port map( A => n5_port, B => n32, Y => n51);
   U87 : XOR2X1 port map( A => N13, B => n73_port, Y => N727);
   U88 : NOR2X1 port map( A => n67, B => n74, Y => n73_port);
   U89 : XOR2X1 port map( A => N9, B => n75, Y => N726);
   U90 : NOR2X1 port map( A => n70, B => n74, Y => n75);
   U91 : XOR2X1 port map( A => N5, B => n76, Y => N725);
   U92 : NOR2X1 port map( A => n62, B => n74, Y => n76);
   U93 : XOR2X1 port map( A => N1, B => n77_port, Y => N724);
   U94 : NOR2X1 port map( A => n30, B => n74, Y => n77_port);
   U95 : NAND3X1 port map( A => n1_port, B => n65_port, C => n52, Y => n74);
   U96 : NOR2X1 port map( A => n11, B => n35, Y => n52);
   U97 : XOR2X1 port map( A => n78, B => n79, Y => n35);
   U98 : XOR2X1 port map( A => n80, B => n81_port, Y => n79);
   U99 : XOR2X1 port map( A => N121, B => N105, Y => n81_port);
   U100 : XOR2X1 port map( A => N89, B => N73, Y => n80);
   U101 : XOR2X1 port map( A => n82, B => n83, Y => n78);
   U102 : XOR2X1 port map( A => n84, B => n85_port, Y => n82);
   U103 : NAND2X1 port map( A => N135, B => N137, Y => n84);
   U104 : XOR2X1 port map( A => n86, B => n87, Y => n32);
   U105 : XOR2X1 port map( A => n88, B => n89_port, Y => n87);
   U106 : XOR2X1 port map( A => N125, B => N109, Y => n89_port);
   U107 : XOR2X1 port map( A => N93, B => N77, Y => n88);
   U108 : XOR2X1 port map( A => n90, B => n91, Y => n86);
   U109 : XOR2X1 port map( A => n92, B => n93_port, Y => n90);
   U110 : NAND2X1 port map( A => N136, B => N137, Y => n92);
   U111 : OAI21X1 port map( A => n45_port, B => n94, C => n95, Y => n65_port);
   U112 : NAND2X1 port map( A => n30, B => n96, Y => n95);
   U113 : OAI21X1 port map( A => n9_port, B => n10, C => n97_port, Y => n96);
   U114 : OAI21X1 port map( A => n21_port, B => n27, C => n62, Y => n97_port);
   U115 : NOR2X1 port map( A => n10, B => n70, Y => n27);
   U116 : NOR2X1 port map( A => n9_port, B => n67, Y => n21_port);
   U117 : NAND2X1 port map( A => n70, B => n67, Y => n94);
   U118 : XOR2X1 port map( A => n98, B => n99, Y => n67);
   U119 : XOR2X1 port map( A => n100, B => n101_port, Y => n99);
   U120 : XOR2X1 port map( A => N29, B => N13, Y => n101_port);
   U121 : XOR2X1 port map( A => N61, B => N45, Y => n100);
   U122 : XOR2X1 port map( A => n102, B => n103, Y => n98);
   U123 : XOR2X1 port map( A => n104, B => n105_port, Y => n102);
   U124 : NAND2X1 port map( A => N132, B => N137, Y => n104);
   U125 : XOR2X1 port map( A => n106, B => n107, Y => n70);
   U126 : XOR2X1 port map( A => n108, B => n109_port, Y => n107);
   U127 : XOR2X1 port map( A => N41, B => N25, Y => n109_port);
   U128 : XOR2X1 port map( A => N9, B => N57, Y => n108);
   U129 : XOR2X1 port map( A => n110, B => n111, Y => n106);
   U130 : XOR2X1 port map( A => n112, B => n113_port, Y => n110);
   U131 : NAND2X1 port map( A => N131, B => N137, Y => n112);
   U132 : NAND2X1 port map( A => n62, B => n7, Y => n45_port);
   U133 : XOR2X1 port map( A => n114, B => n115, Y => n62);
   U134 : XOR2X1 port map( A => n116, B => n117_port, Y => n115);
   U135 : XOR2X1 port map( A => N37, B => N21, Y => n117_port);
   U136 : XOR2X1 port map( A => N53, B => N5, Y => n116);
   U137 : XOR2X1 port map( A => n118, B => n111, Y => n114);
   U138 : XNOR2X1 port map( A => n119, B => n120, Y => n111);
   U139 : XOR2X1 port map( A => N97, B => N109, Y => n120);
   U140 : XNOR2X1 port map( A => N101, B => N105, Y => n119);
   U141 : XOR2X1 port map( A => n121_port, B => n103, Y => n118);
   U142 : XNOR2X1 port map( A => n122, B => n123, Y => n103);
   U143 : XOR2X1 port map( A => N125, B => N121, Y => n123);
   U144 : XOR2X1 port map( A => N113, B => n15, Y => n122);
   U145 : NAND2X1 port map( A => N130, B => N137, Y => n121_port);
   U146 : NAND2X1 port map( A => n37_port, B => n3, Y => n46);
   U147 : XOR2X1 port map( A => n124, B => n125_port, Y => n39);
   U148 : XOR2X1 port map( A => n126, B => n127, Y => n125_port);
   U149 : XOR2X1 port map( A => N65, B => N113, Y => n127);
   U150 : XOR2X1 port map( A => N97, B => N81, Y => n126);
   U151 : XOR2X1 port map( A => n128, B => n85_port, Y => n124);
   U152 : XNOR2X1 port map( A => n129_port, B => n130_port, Y => n85_port);
   U153 : XOR2X1 port map( A => N9, B => N5, Y => n130_port);
   U154 : XNOR2X1 port map( A => N1, B => N13, Y => n129_port);
   U155 : XOR2X1 port map( A => n131_port, B => n93_port, Y => n128);
   U156 : XNOR2X1 port map( A => n132_port, B => n133_port, Y => n93_port);
   U157 : XOR2X1 port map( A => N29, B => N25, Y => n133_port);
   U158 : XNOR2X1 port map( A => N17, B => N21, Y => n132_port);
   U159 : NAND2X1 port map( A => N133, B => N137, Y => n131_port);
   U160 : XOR2X1 port map( A => n134_port, B => n135_port, Y => n37_port);
   U161 : XOR2X1 port map( A => n136_port, B => n137_port, Y => n135_port);
   U162 : XOR2X1 port map( A => N117, B => N101, Y => n137_port);
   U163 : XOR2X1 port map( A => N85, B => N69, Y => n136_port);
   U164 : XOR2X1 port map( A => n138, B => n83, Y => n134_port);
   U165 : XNOR2X1 port map( A => n139, B => n140, Y => n83);
   U166 : XOR2X1 port map( A => N45, B => N41, Y => n140);
   U167 : XNOR2X1 port map( A => N33, B => N37, Y => n139);
   U168 : XOR2X1 port map( A => n141, B => n91, Y => n138);
   U169 : XNOR2X1 port map( A => n142, B => n143, Y => n91);
   U170 : XOR2X1 port map( A => N61, B => N57, Y => n143);
   U171 : XOR2X1 port map( A => n13_port, B => N53, Y => n142);
   U172 : NAND2X1 port map( A => N137, B => N134, Y => n141);
   U173 : XOR2X1 port map( A => n144, B => n145, Y => n30);
   U174 : XOR2X1 port map( A => n146, B => n147, Y => n145);
   U175 : XOR2X1 port map( A => N17, B => N1, Y => n147);
   U176 : XOR2X1 port map( A => N49, B => N33, Y => n146);
   U177 : XOR2X1 port map( A => n148, B => n113_port, Y => n144);
   U178 : XNOR2X1 port map( A => n149, B => n150, Y => n113_port);
   U179 : XOR2X1 port map( A => N77, B => N73, Y => n150);
   U180 : XOR2X1 port map( A => n14, B => N69, Y => n149);
   U181 : XOR2X1 port map( A => n151, B => n105_port, Y => n148);
   U182 : XNOR2X1 port map( A => n152, B => n153, Y => n105_port);
   U183 : XOR2X1 port map( A => N93, B => N89, Y => n153);
   U184 : XNOR2X1 port map( A => N81, B => N85, Y => n152);
   U185 : NAND2X1 port map( A => N129, B => N137, Y => n151);

end SYN_verilog;

library IEEE;

use IEEE.std_logic_1164.all;

entity c499_clk_opFF is

   port( clk, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53
         , N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, 
         N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135
         , N136, N137 : in std_logic;  Qout_N724, Qout_N725, Qout_N726, 
         Qout_N727, Qout_N728, Qout_N729, Qout_N730, Qout_N731, Qout_N732, 
         Qout_N733, Qout_N734, Qout_N735, Qout_N736, Qout_N737, Qout_N738, 
         Qout_N739, Qout_N740, Qout_N741, Qout_N742, Qout_N743, Qout_N744, 
         Qout_N745, Qout_N746, Qout_N747, Qout_N748, Qout_N749, Qout_N750, 
         Qout_N751, Qout_N752, Qout_N753, Qout_N754, Qout_N755 : out std_logic
         );

end c499_clk_opFF;

architecture SYN_verilog of c499_clk_opFF is

   component dff_0
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_1
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_2
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_3
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_4
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_5
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_6
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_7
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_8
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_9
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_10
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_11
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_12
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_13
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_14
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_15
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_16
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_17
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_18
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_19
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_20
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_21
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_22
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_23
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_24
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_25
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_26
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_27
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_28
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_29
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_30
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_31
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_32
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_33
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_34
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_35
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_36
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_37
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_38
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_39
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_40
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_41
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_42
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_43
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_44
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_45
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_46
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_47
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_48
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_49
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_50
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_51
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_52
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_53
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_54
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_55
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_56
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_57
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_58
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_59
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_60
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_61
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_62
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_63
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_64
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_65
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_66
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_67
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_68
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_69
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_70
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_71
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_72
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_73
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_74
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_75
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_76
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_77
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_78
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_79
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_80
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_81
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_82
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_83
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_84
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_85
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_86
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_87
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_88
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_89
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_90
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_91
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_92
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_93
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_94
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_95
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_96
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_97
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_98
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_99
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_100
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_101
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_102
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_103
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component dff_104
      port( q : out std_logic;  d, clk : in std_logic);
   end component;
   
   component c499
      port( N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, 
            N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, 
            N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, 
            N135, N136, N137 : in std_logic;  N724, N725, N726, N727, N728, 
            N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, 
            N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, 
            N751, N752, N753, N754, N755 : out std_logic);
   end component;
   
   signal IN_N1, IN_N5, IN_N9, IN_N13, IN_N17, IN_N21, IN_N25, IN_N29, IN_N33, 
      IN_N37, IN_N41, IN_N45, IN_N49, IN_N53, IN_N57, IN_N61, IN_N65, IN_N69, 
      IN_N73, IN_N77, IN_N81, IN_N85, IN_N89, IN_N93, IN_N97, IN_N101, IN_N105,
      IN_N109, IN_N113, IN_N117, IN_N121, IN_N125, IN_N129, IN_N130, IN_N131, 
      IN_N132, IN_N133, IN_N134, IN_N135, IN_N136, IN_N137, N724, N725, N726, 
      N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, 
      N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, 
      N751, N752, N753, N754, N755, Q_N724, Q_N725, Q_N726, Q_N727, Q_N728, 
      Q_N729, Q_N730, Q_N731, Q_N732, Q_N733, Q_N734, Q_N735, Q_N736, Q_N737, 
      Q_N738, Q_N739, Q_N740, Q_N741, Q_N742, Q_N743, Q_N744, Q_N745, Q_N746, 
      Q_N747, Q_N748, Q_N749, Q_N750, Q_N751, Q_N752, Q_N753, Q_N754, Q_N755 : 
      std_logic;

begin
   
   c0 : c499 port map( N1 => IN_N1, N5 => IN_N5, N9 => IN_N9, N13 => IN_N13, 
                           N17 => IN_N17, N21 => IN_N21, N25 => IN_N25, N29 => 
                           IN_N29, N33 => IN_N33, N37 => IN_N37, N41 => IN_N41,
                           N45 => IN_N45, N49 => IN_N49, N53 => IN_N53, N57 => 
                           IN_N57, N61 => IN_N61, N65 => IN_N65, N69 => IN_N69,
                           N73 => IN_N73, N77 => IN_N77, N81 => IN_N81, N85 => 
                           IN_N85, N89 => IN_N89, N93 => IN_N93, N97 => IN_N97,
                           N101 => IN_N101, N105 => IN_N105, N109 => IN_N109, 
                           N113 => IN_N113, N117 => IN_N117, N121 => IN_N121, 
                           N125 => IN_N125, N129 => IN_N129, N130 => IN_N130, 
                           N131 => IN_N131, N132 => IN_N132, N133 => IN_N133, 
                           N134 => IN_N134, N135 => IN_N135, N136 => IN_N136, 
                           N137 => IN_N137, N724 => N724, N725 => N725, N726 =>
                           N726, N727 => N727, N728 => N728, N729 => N729, N730
                           => N730, N731 => N731, N732 => N732, N733 => N733, 
                           N734 => N734, N735 => N735, N736 => N736, N737 => 
                           N737, N738 => N738, N739 => N739, N740 => N740, N741
                           => N741, N742 => N742, N743 => N743, N744 => N744, 
                           N745 => N745, N746 => N746, N747 => N747, N748 => 
                           N748, N749 => N749, N750 => N750, N751 => N751, N752
                           => N752, N753 => N753, N754 => N754, N755 => N755);
   iDFF_1 : dff_104 port map( q => IN_N1, d => N1, clk => clk);
   iDFF_2 : dff_103 port map( q => IN_N5, d => N5, clk => clk);
   iDFF_3 : dff_102 port map( q => IN_N9, d => N9, clk => clk);
   iDFF_4 : dff_101 port map( q => IN_N13, d => N13, clk => clk);
   iDFF_5 : dff_100 port map( q => IN_N17, d => N17, clk => clk);
   iDFF_6 : dff_99 port map( q => IN_N21, d => N21, clk => clk);
   iDFF_7 : dff_98 port map( q => IN_N25, d => N25, clk => clk);
   iDFF_8 : dff_97 port map( q => IN_N29, d => N29, clk => clk);
   iDFF_9 : dff_96 port map( q => IN_N33, d => N33, clk => clk);
   iDFF_10 : dff_95 port map( q => IN_N37, d => N37, clk => clk);
   iDFF_11 : dff_94 port map( q => IN_N41, d => N41, clk => clk);
   iDFF_12 : dff_93 port map( q => IN_N45, d => N45, clk => clk);
   iDFF_13 : dff_92 port map( q => IN_N49, d => N49, clk => clk);
   iDFF_14 : dff_91 port map( q => IN_N53, d => N53, clk => clk);
   iDFF_15 : dff_90 port map( q => IN_N57, d => N57, clk => clk);
   iDFF_16 : dff_89 port map( q => IN_N61, d => N61, clk => clk);
   iDFF_17 : dff_88 port map( q => IN_N65, d => N65, clk => clk);
   iDFF_18 : dff_87 port map( q => IN_N69, d => N69, clk => clk);
   iDFF_19 : dff_86 port map( q => IN_N73, d => N73, clk => clk);
   iDFF_20 : dff_85 port map( q => IN_N77, d => N77, clk => clk);
   iDFF_21 : dff_84 port map( q => IN_N81, d => N81, clk => clk);
   iDFF_22 : dff_83 port map( q => IN_N85, d => N85, clk => clk);
   iDFF_23 : dff_82 port map( q => IN_N89, d => N89, clk => clk);
   iDFF_24 : dff_81 port map( q => IN_N93, d => N93, clk => clk);
   iDFF_25 : dff_80 port map( q => IN_N97, d => N97, clk => clk);
   iDFF_26 : dff_79 port map( q => IN_N101, d => N101, clk => clk);
   iDFF_27 : dff_78 port map( q => IN_N105, d => N105, clk => clk);
   iDFF_28 : dff_77 port map( q => IN_N109, d => N109, clk => clk);
   iDFF_29 : dff_76 port map( q => IN_N113, d => N113, clk => clk);
   iDFF_30 : dff_75 port map( q => IN_N117, d => N117, clk => clk);
   iDFF_31 : dff_74 port map( q => IN_N121, d => N121, clk => clk);
   iDFF_32 : dff_73 port map( q => IN_N125, d => N125, clk => clk);
   iDFF_33 : dff_72 port map( q => IN_N129, d => N129, clk => clk);
   iDFF_34 : dff_71 port map( q => IN_N130, d => N130, clk => clk);
   iDFF_35 : dff_70 port map( q => IN_N131, d => N131, clk => clk);
   iDFF_36 : dff_69 port map( q => IN_N132, d => N132, clk => clk);
   iDFF_37 : dff_68 port map( q => IN_N133, d => N133, clk => clk);
   iDFF_38 : dff_67 port map( q => IN_N134, d => N134, clk => clk);
   iDFF_39 : dff_66 port map( q => IN_N135, d => N135, clk => clk);
   iDFF_40 : dff_65 port map( q => IN_N136, d => N136, clk => clk);
   iDFF_41 : dff_64 port map( q => IN_N137, d => N137, clk => clk);
   DFF_1_inst : dff_63 port map( q => Q_N724, d => N724, clk => clk);
   DFF_2_inst : dff_62 port map( q => Q_N725, d => N725, clk => clk);
   DFF_3_inst : dff_61 port map( q => Q_N726, d => N726, clk => clk);
   DFF_4_inst : dff_60 port map( q => Q_N727, d => N727, clk => clk);
   DFF_5_inst : dff_59 port map( q => Q_N728, d => N728, clk => clk);
   DFF_6_inst : dff_58 port map( q => Q_N729, d => N729, clk => clk);
   DFF_7_inst : dff_57 port map( q => Q_N730, d => N730, clk => clk);
   DFF_8_inst : dff_56 port map( q => Q_N731, d => N731, clk => clk);
   DFF_9_inst : dff_55 port map( q => Q_N732, d => N732, clk => clk);
   DFF_10_inst : dff_54 port map( q => Q_N733, d => N733, clk => clk);
   DFF_11_inst : dff_53 port map( q => Q_N734, d => N734, clk => clk);
   DFF_12_inst : dff_52 port map( q => Q_N735, d => N735, clk => clk);
   DFF_13_inst : dff_51 port map( q => Q_N736, d => N736, clk => clk);
   DFF_14_inst : dff_50 port map( q => Q_N737, d => N737, clk => clk);
   DFF_15_inst : dff_49 port map( q => Q_N738, d => N738, clk => clk);
   DFF_16_inst : dff_48 port map( q => Q_N739, d => N739, clk => clk);
   DFF_17_inst : dff_47 port map( q => Q_N740, d => N740, clk => clk);
   DFF_18_inst : dff_46 port map( q => Q_N741, d => N741, clk => clk);
   DFF_19_inst : dff_45 port map( q => Q_N742, d => N742, clk => clk);
   DFF_20_inst : dff_44 port map( q => Q_N743, d => N743, clk => clk);
   DFF_21_inst : dff_43 port map( q => Q_N744, d => N744, clk => clk);
   DFF_22_inst : dff_42 port map( q => Q_N745, d => N745, clk => clk);
   DFF_23_inst : dff_41 port map( q => Q_N746, d => N746, clk => clk);
   DFF_24_inst : dff_40 port map( q => Q_N747, d => N747, clk => clk);
   DFF_25_inst : dff_39 port map( q => Q_N748, d => N748, clk => clk);
   DFF_26_inst : dff_38 port map( q => Q_N749, d => N749, clk => clk);
   DFF_27_inst : dff_37 port map( q => Q_N750, d => N750, clk => clk);
   DFF_28_inst : dff_36 port map( q => Q_N751, d => N751, clk => clk);
   DFF_29_inst : dff_35 port map( q => Q_N752, d => N752, clk => clk);
   DFF_30_inst : dff_34 port map( q => Q_N753, d => N753, clk => clk);
   DFF_31_inst : dff_33 port map( q => Q_N754, d => N754, clk => clk);
   DFF_32_inst : dff_32 port map( q => Q_N755, d => N755, clk => clk);
   oDFF_1 : dff_31 port map( q => Qout_N724, d => Q_N724, clk => clk);
   oDFF_2 : dff_30 port map( q => Qout_N725, d => Q_N725, clk => clk);
   oDFF_3 : dff_29 port map( q => Qout_N726, d => Q_N726, clk => clk);
   oDFF_4 : dff_28 port map( q => Qout_N727, d => Q_N727, clk => clk);
   oDFF_5 : dff_27 port map( q => Qout_N728, d => Q_N728, clk => clk);
   oDFF_6 : dff_26 port map( q => Qout_N729, d => Q_N729, clk => clk);
   oDFF_7 : dff_25 port map( q => Qout_N730, d => Q_N730, clk => clk);
   oDFF_8 : dff_24 port map( q => Qout_N731, d => Q_N731, clk => clk);
   oDFF_9 : dff_23 port map( q => Qout_N732, d => Q_N732, clk => clk);
   oDFF_10 : dff_22 port map( q => Qout_N733, d => Q_N733, clk => clk);
   oDFF_11 : dff_21 port map( q => Qout_N734, d => Q_N734, clk => clk);
   oDFF_12 : dff_20 port map( q => Qout_N735, d => Q_N735, clk => clk);
   oDFF_13 : dff_19 port map( q => Qout_N736, d => Q_N736, clk => clk);
   oDFF_14 : dff_18 port map( q => Qout_N737, d => Q_N737, clk => clk);
   oDFF_15 : dff_17 port map( q => Qout_N738, d => Q_N738, clk => clk);
   oDFF_16 : dff_16 port map( q => Qout_N739, d => Q_N739, clk => clk);
   oDFF_17 : dff_15 port map( q => Qout_N740, d => Q_N740, clk => clk);
   oDFF_18 : dff_14 port map( q => Qout_N741, d => Q_N741, clk => clk);
   oDFF_19 : dff_13 port map( q => Qout_N742, d => Q_N742, clk => clk);
   oDFF_20 : dff_12 port map( q => Qout_N743, d => Q_N743, clk => clk);
   oDFF_21 : dff_11 port map( q => Qout_N744, d => Q_N744, clk => clk);
   oDFF_22 : dff_10 port map( q => Qout_N745, d => Q_N745, clk => clk);
   oDFF_23 : dff_9 port map( q => Qout_N746, d => Q_N746, clk => clk);
   oDFF_24 : dff_8 port map( q => Qout_N747, d => Q_N747, clk => clk);
   oDFF_25 : dff_7 port map( q => Qout_N748, d => Q_N748, clk => clk);
   oDFF_26 : dff_6 port map( q => Qout_N749, d => Q_N749, clk => clk);
   oDFF_27 : dff_5 port map( q => Qout_N750, d => Q_N750, clk => clk);
   oDFF_28 : dff_4 port map( q => Qout_N751, d => Q_N751, clk => clk);
   oDFF_29 : dff_3 port map( q => Qout_N752, d => Q_N752, clk => clk);
   oDFF_30 : dff_2 port map( q => Qout_N753, d => Q_N753, clk => clk);
   oDFF_31 : dff_1 port map( q => Qout_N754, d => Q_N754, clk => clk);
   oDFF_32 : dff_0 port map( q => Qout_N755, d => Q_N755, clk => clk);

end SYN_verilog;
