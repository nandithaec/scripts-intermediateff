library verilog;
use verilog.vl_types.all;
entity XOR2X1 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        Y               : out    vl_logic
    );
end XOR2X1;
