library verilog;
use verilog.vl_types.all;
entity AOI21X1 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        Y               : out    vl_logic
    );
end AOI21X1;
