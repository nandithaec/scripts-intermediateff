****Template spice file***

.include ../glitch_osu018_stdcells_correct_vdd_gnd.sp
**.include /cad/digital/rtl2gds/rtl2gds_install/LIB/lib/tsmc018/lib/tsmc018.m
.include ../tsmc018.m

**********Subckt begins*********

.SUBCKT c499_clk_opFF
+       clk N1 N5 N9 N13 N17 N21 N25 N29 N33 N37 N41 N45 N49 N53 N57 N61 N65 N69
+       N73 N77 N81 N85 N89 N93 N97 N101 N105 N109 N113 N117 N121 N125 N129 N130
+       N131 N132 N133 N134 N135 N136 N137 Qout_N724 Qout_N725 Qout_N726
+       Qout_N727 Qout_N728 Qout_N729 Qout_N730 Qout_N731 Qout_N732 Qout_N733
+       Qout_N734 Qout_N735 Qout_N736 Qout_N737 Qout_N738 Qout_N739 Qout_N740
+       Qout_N741 Qout_N742 Qout_N743 Qout_N744 Qout_N745 Qout_N746 Qout_N747
+       Qout_N748 Qout_N749 Qout_N750 Qout_N751 Qout_N752 Qout_N753 Qout_N754
+       Qout_N755
C1 iDFF_4_q_reg:D 0 1.86274e-16
C2 N13 0 4.18369e-15
C3 N13:4 0 1.65296e-15
R1 iDFF_4_q_reg:D N13:4 12.3333
R2 N13 N13:4 16.3833
C4 N1 0 3.52533e-15
C5 iDFF_1_q_reg:D 0 1.1313e-16
C6 N1:2 0 1.03808e-15
R3 N1 N1:2 43.05
R4 iDFF_1_q_reg:D N1:2 10.7333
C7 N131 0 4.77275e-15
C8 iDFF_35_q_reg:D 0 1.47374e-16
R5 N131 iDFF_35_q_reg:D 24.5167
C9 Qout_N728 0 2.59069e-15
C10 oDFF_5_q_reg:Q 0 1.04278e-16
R6 oDFF_5_q_reg:Q Qout_N728 20.1833
C11 Qout_N739 0 5.96796e-17
C12 oDFF_16_q_reg:Q 0 3.26358e-15
R7 oDFF_16_q_reg:Q Qout_N739 23.5167
C13 DFF_4_q_reg:D 0 8.8421e-16
C14 c0_U87:Y 0 1.18219e-16
C15 N727:2 0 7.70145e-16
R8 c0_U87:Y N727:2 24.2667
R9 DFF_4_q_reg:D N727:2 9.26667
C16 oDFF_4_q_reg:D 0 6.51495e-16
C17 DFF_4_q_reg:Q 0 1.35551e-15
R10 DFF_4_q_reg:Q oDFF_4_q_reg:D 20.1333
C18 oDFF_6_q_reg:Q 0 4.97621e-16
C19 Qout_N729 0 3.53716e-15
C20 Qout_N729:5 0 9.1377e-16
R11 oDFF_6_q_reg:Q Qout_N729:5 44.3067
R12 Qout_N729 Qout_N729:5 16.3
C21 N5 0 2.6236e-15
C22 iDFF_2_q_reg:D 0 5.12382e-16
C23 N5:3 0 1.84488e-15
R13 N5 N5:3 12.8333
R14 iDFF_2_q_reg:D N5:3 44.5733
C24 N9 0 2.11658e-15
C25 iDFF_3_q_reg:D 0 1.8127e-16
C26 N9:3 0 1.35559e-15
R15 N9 N9:3 18.7883
R16 iDFF_3_q_reg:D N9:3 18.2
C27 N25 0 2.83509e-15
C28 iDFF_7_q_reg:D 0 1.51453e-16
R17 N25 iDFF_7_q_reg:D 27.2333
C29 Qout_N725 0 1.30489e-15
C30 oDFF_2_q_reg:Q 0 2.05038e-15
R18 oDFF_2_q_reg:Q Qout_N725 26.7
C31 Qout_N730 0 1.25546e-15
C32 oDFF_7_q_reg:Q 0 1.97271e-15
R19 oDFF_7_q_reg:Q Qout_N730 26.1667
C33 Qout_N731 0 1.5057e-15
C34 oDFF_8_q_reg:Q 0 2.471e-15
R20 oDFF_8_q_reg:Q Qout_N731 29.1
C35 c0_U88:A 0 7.43027e-16
C36 c0_U118:Y 0 6.13781e-16
C37 c0_U10:A 0 3.23184e-16
C38 c0_U117:B 0 1.97746e-16
C39 c0_U116:B 0 1.25679e-16
C40 c0_U78:A 0 1.40273e-16
C41 c0_n67:10 0 1.52049e-15
C42 c0_n67:12 0 1.38684e-15
C43 c0_n67:14 0 1.23322e-15
R21 c0_U88:A c0_n67:10 10.4
R22 c0_U118:Y c0_n67:10 23.2
R23 c0_U118:Y c0_n67:12 14.0667
R24 c0_U116:B c0_U10:A 52.7735
R25 c0_U10:A c0_n67:14 37.585
R26 c0_U117:B c0_n67:14 22.7333
R27 c0_U116:B c0_n67:14 31.5776
R28 c0_U78:A c0_n67:10 7.66667
R29 c0_n67:12 c0_n67:14 17.0667
C44 iDFF_2_q_reg:Q 0 1.07223e-15
C45 c0_U153:B 0 2.80526e-16
C46 c0_U136:B 0 6.93381e-16
C47 c0_U91:A 0 9.29894e-16
C48 IN_N5:5 0 1.72925e-15
R30 iDFF_2_q_reg:Q IN_N5:5 11.7333
R31 iDFF_2_q_reg:Q c0_U136:B 29.8667
R32 c0_U91:A IN_N5:5 22.2667
R33 c0_U136:B c0_U153:B 1.06667
C49 iDFF_3_q_reg:Q 0 1.05656e-15
C50 c0_U153:A 0 3.5829e-16
C51 c0_U128:A 0 7.40645e-16
C52 c0_U89:A 0 4.46112e-16
R34 iDFF_3_q_reg:Q c0_U89:A 15.4667
R35 c0_U89:A c0_U128:A 1.33333
R36 c0_U128:A c0_U153:A 28.2667
C53 iDFF_4_q_reg:Q 0 3.38649e-16
C54 c0_U154:B 0 8.16303e-16
C55 c0_U120:B 0 1.81086e-16
C56 c0_U87:A 0 9.09717e-17
C57 IN_N13:4 0 1.39896e-15
R37 iDFF_4_q_reg:Q c0_U87:A 0.266667
R38 iDFF_4_q_reg:Q IN_N13:4 20.7333
R39 c0_U120:B c0_U154:B 15.4
R40 c0_U154:B IN_N13:4 11.4
C58 iDFF_5_q_reg:Q 0 5.17452e-16
C59 c0_U175:A 0 5.17831e-16
C60 c0_U158:A 0 1.79475e-16
C61 c0_U83:A 0 7.57042e-16
C62 IN_N17:6 0 1.45672e-15
R41 iDFF_5_q_reg:Q IN_N17:6 222.721
R42 iDFF_5_q_reg:Q c0_U175:A 94.1903
R43 iDFF_5_q_reg:Q c0_U83:A 35.9402
R44 c0_U83:A IN_N17:6 222.721
R45 c0_U83:A c0_U175:A 94.1903
R46 c0_U158:A IN_N17:6 9.73333
R47 c0_U175:A IN_N17:6 24.9198
C63 iDFF_7_q_reg:Q 0 1.0252e-15
C64 c0_U157:B 0 1.31522e-15
C65 c0_U127:B 0 5.75038e-16
C66 c0_U79:A 0 6.58727e-16
R48 iDFF_7_q_reg:Q c0_U79:A 66.9325
R49 iDFF_7_q_reg:Q c0_U127:B 91.3349
R50 iDFF_7_q_reg:Q c0_U157:B 54.8562
R51 c0_U79:A c0_U127:B 18.6935
R52 c0_U79:A c0_U157:B 67.4902
R53 c0_U127:B c0_U157:B 92.0961
C67 iDFF_8_q_reg:Q 0 5.15208e-16
C68 c0_U157:A 0 1.17577e-15
C69 c0_U120:A 0 3.00947e-16
C70 c0_U77:A 0 7.73351e-16
R54 iDFF_8_q_reg:Q c0_U157:A 28.8667
R55 c0_U77:A c0_U157:A 55.3531
R56 c0_U77:A c0_U120:A 18.9181
R57 c0_U120:A c0_U157:A 45.6346
C71 iDFF_11_q_reg:Q 0 1.00342e-15
C72 c0_U166:B 0 4.11668e-16
C73 c0_U127:A 0 3.01238e-16
C74 c0_U69:A 0 1.98829e-16
C75 IN_N41:5 0 2.51286e-15
R58 iDFF_11_q_reg:Q IN_N41:5 15.6667
R59 iDFF_11_q_reg:Q c0_U69:A 20.7867
R60 iDFF_11_q_reg:Q c0_U166:B 51.9667
R61 c0_U69:A c0_U166:B 1.91582
R62 c0_U127:A IN_N41:5 21.1333
C76 DFF_2_q_reg:D 0 2.68985e-15
C77 c0_U91:Y 0 5.47628e-16
R63 c0_U91:Y DFF_2_q_reg:D 48.1333
C78 DFF_3_q_reg:D 0 5.421e-16
C79 c0_U89:Y 0 5.6546e-16
R64 c0_U89:Y DFF_3_q_reg:D 28.5333
C80 DFF_7_q_reg:D 0 1.09851e-16
C81 c0_U79:Y 0 1.50949e-16
C82 N730:2 0 9.94327e-16
R65 c0_U79:Y N730:2 21.3333
R66 DFF_7_q_reg:D N730:2 6.73333
C83 DFF_8_q_reg:D 0 7.73615e-16
C84 c0_U77:Y 0 4.36565e-16
R67 c0_U77:Y DFF_8_q_reg:D 31.1333
C85 oDFF_2_q_reg:D 0 7.15313e-16
C86 DFF_2_q_reg:Q 0 4.55699e-16
R68 DFF_2_q_reg:Q oDFF_2_q_reg:D 28.4
C87 c0_U171:A 0 9.12304e-16
C88 c0_U64:A 0 1.30447e-16
C89 c0_U13:Y 0 1.52357e-16
C90 c0_n13:3 0 2.89127e-15
R69 c0_U13:Y c0_n13:3 14.9333
R70 c0_U64:A c0_n13:3 18.8
R71 c0_U171:A c0_n13:3 16.1333
C91 c0_U77:B 0 2.06585e-16
R72 c0_U78:Y c0_U77:B 0.533333
C92 c0_U79:B 0 1.91307e-16
R73 c0_U80:Y c0_U79:B 0.533333
C93 c0_U84:Y 0 3.93614e-16
C94 c0_U83:B 0 9.65694e-16
R74 c0_U84:Y c0_U83:B 28.8667
C95 c0_U88:Y 0 4.66945e-16
C96 c0_U87:B 0 6.08424e-16
R75 c0_U88:Y c0_U87:B 16.4
C97 c0_U90:Y 0 4.84601e-16
C98 c0_U89:B 0 7.83641e-16
R76 c0_U90:Y c0_U89:B 30.4667
C99 c0_U92:Y 0 1.17899e-16
C100 c0_U91:B 0 9.44674e-16
C101 c0_n76:3 0 1.31496e-15
R77 c0_U92:Y c0_n76:3 9.73333
R78 c0_U91:B c0_n76:3 22.2
C102 c0_U94:Y 0 3.72964e-16
C103 c0_U93:B 0 1.94042e-15
R79 c0_U94:Y c0_U93:B 21
C104 c0_U113:Y 0 8.4425e-16
C105 c0_U112:B 0 1.16093e-16
R80 c0_U113:Y c0_U112:B 3.53333
C106 c0_U119:Y 0 3.99178e-16
C107 c0_U118:B 0 5.40751e-16
R81 c0_U119:Y c0_U118:B 28.6
C108 c0_U120:Y 0 5.19484e-16
C109 c0_U119:B 0 2.4519e-16
C110 c0_n101:2 0 1.03915e-15
R82 c0_U120:Y c0_n101:2 8.06667
R83 c0_U119:B c0_n101:2 21.0667
C111 c0_U128:Y 0 3.53239e-16
C112 c0_U126:A 0 9.57927e-16
R84 c0_U128:Y c0_U126:A 29.6
C113 c0_U127:Y 0 8.40905e-16
C114 c0_U126:B 0 7.91937e-16
R85 c0_U127:Y c0_U126:B 30.9333
C115 c0_U154:Y 0 4.66181e-16
C116 c0_U152:A 0 6.66149e-16
C117 c0_n129:2 0 8.07861e-16
R86 c0_U154:Y c0_n129:2 14.8667
R87 c0_U152:A c0_n129:2 30.6
C118 c0_U158:Y 0 5.59755e-16
C119 c0_U156:A 0 1.57943e-16
R88 c0_U158:Y c0_U156:A 14.4667
C120 c0_U157:Y 0 1.85122e-15
C121 c0_U156:B 0 2.21411e-16
C122 c0_n133:2 0 2.65116e-15
R89 c0_U157:Y c0_n133:2 19.2667
R90 c0_U156:B c0_n133:2 18.6667
C123 c0_U171:Y 0 1.32662e-16
C124 c0_U169:A 0 6.72149e-16
R91 c0_U171:Y c0_U169:A 15.2667
C125 c0_U170:Y 0 5.49239e-16
C126 c0_U169:B 0 1.28559e-16
R92 c0_U170:Y c0_U169:B 2.2
C127 c0_U174:Y 0 1.49705e-16
C128 c0_U173:B 0 1.39723e-16
C129 c0_n145:2 0 9.75803e-16
R93 c0_U174:Y c0_n145:2 20.2667
R94 c0_U173:B c0_n145:2 9.06667
C130 c0_U175:Y 0 1.01111e-15
C131 c0_U174:B 0 3.98766e-16
R95 c0_U175:Y c0_U174:B 29.4
C132 c0_U80:A 0 5.59786e-16
C133 c0_U125:Y 0 5.039e-16
C134 c0_U90:A 0 3.05742e-16
C135 c0_U9:A 0 7.46529e-17
C136 c0_U117:A 0 5.9768e-16
C137 c0_U115:B 0 4.98343e-16
C138 c0_n70:8 0 9.76542e-16
C139 c0_n70:10 0 5.50039e-16
R96 c0_U80:A c0_n70:8 8.06667
R97 c0_U125:Y c0_U117:A 15.4667
R98 c0_U90:A c0_n70:8 154.158
R99 c0_U90:A c0_n70:10 17.4818
R100 c0_U9:A c0_n70:10 13.1333
R101 c0_U117:A c0_U115:B 28.8333
R102 c0_U117:A c0_n70:10 27.2606
R103 c0_U115:B c0_n70:10 34.6
R104 c0_n70:8 c0_n70:10 34.6068
C140 iDFF_12_q_reg:Q 0 1.08802e-15
C141 c0_U166:A 0 6.4052e-16
C142 c0_U121:B 0 1.14035e-16
C143 c0_U67:A 0 4.13073e-16
C144 IN_N45:6 0 2.48068e-15
R105 iDFF_12_q_reg:Q IN_N45:6 61.3045
R106 iDFF_12_q_reg:Q c0_U67:A 41.8335
R107 c0_U67:A IN_N45:6 54.5208
R108 c0_U121:B IN_N45:6 12.8
R109 c0_U166:A IN_N45:6 17.2667
C145 DFF_6_q_reg:D 0 1.01483e-15
C146 c0_U81:Y 0 2.03173e-16
R110 c0_U81:Y DFF_6_q_reg:D 27.7333
C147 DFF_11_q_reg:D 0 7.16478e-16
C148 c0_U69:Y 0 5.40325e-16
R111 c0_U69:Y DFF_11_q_reg:D 28.2667
C149 oDFF_11_q_reg:D 0 5.60102e-16
C150 DFF_11_q_reg:Q 0 6.706e-16
R112 DFF_11_q_reg:Q oDFF_11_q_reg:D 29.2
C151 c0_U70:Y 0 2.09284e-16
C152 c0_U69:B 0 1.38772e-16
C153 c0_n60:2 0 1.80932e-15
R113 c0_U70:Y c0_n60:2 27.5333
R114 c0_U69:B c0_n60:2 7.06667
C154 c0_U121:Y 0 9.31027e-17
C155 c0_U119:A 0 1.49559e-15
C156 c0_n100:3 0 8.84166e-16
C157 c0_n100:4 0 1.28258e-15
R115 c0_U121:Y c0_n100:4 10.7333
R116 c0_U119:A c0_n100:3 11.7333
R117 c0_n100:3 c0_n100:4 33.2667
C158 c0_U129:Y 0 1.65313e-16
C159 c0_U125:A 0 2.02963e-16
C160 c0_n106:2 0 1.78562e-15
R118 c0_U129:Y c0_n106:2 24
R119 c0_U125:A c0_n106:2 7.06667
C161 c0_U126:Y 0 1.77026e-15
C162 c0_U125:B 0 3.84733e-16
R120 c0_U126:Y c0_U125:B 30.5333
C163 c0_U137:Y 0 1.55944e-16
C164 c0_U133:A 0 8.77768e-16
C165 c0_n114:2 0 1.72454e-15
R121 c0_U137:Y c0_n114:2 24
R122 c0_U133:A c0_n114:2 9.26667
C166 c0_U134:Y 0 5.57517e-16
C167 c0_U133:B 0 8.4436e-16
R123 c0_U134:Y c0_U133:B 29.3333
C168 c0_U136:Y 0 1.31868e-15
C169 c0_U134:A 0 4.28184e-16
R124 c0_U136:Y c0_U134:A 29.4667
C170 c0_U135:Y 0 4.24917e-16
C171 c0_U134:B 0 2.2872e-16
R125 c0_U135:Y c0_U134:B 1.93333
C172 c0_U153:Y 0 9.41848e-17
C173 c0_U152:B 0 1.30198e-15
C174 c0_n130:5 0 1.25687e-15
R126 c0_U153:Y c0_n130:5 8.06667
R127 c0_U152:B c0_n130:5 24.1333
C175 c0_U170:B 0 2.36352e-16
C176 iDFF_15_q_reg:Q 0 4.62419e-16
C177 c0_U128:B 0 6.5553e-16
C178 iDFF_15_q_reg:Q 0 7.56606e-16
C179 c0_U60:A 0 5.76794e-16
C180 IN_N57:7 0 2.81047e-15
R128 c0_U170:B IN_N57:7 24.3333
R129 iDFF_15_q_reg:Q c0_U128:B 29.6667
R130 iDFF_15_q_reg:Q IN_N57:7 9.66667
R131 c0_U60:A IN_N57:7 26.0667
C181 c0_U61:B 0 6.45132e-16
C182 c0_U113:A 0 5.47795e-16
C183 c0_U70:B 0 2.3014e-16
C184 c0_U116:A 0 1.23087e-16
C185 c0_U9:Y 0 3.529e-16
C186 c0_n9:11 0 2.02771e-15
R132 c0_U70:B c0_U61:B 56.5543
R133 c0_U61:B c0_n9:11 61.8562
R134 c0_U113:A c0_n9:11 22.2
R135 c0_U70:B c0_n9:11 15.1099
R136 c0_U116:A c0_U9:Y 1.33333
R137 c0_U116:A c0_n9:11 7.06667
C187 c0_U115:A 0 1.39705e-16
C188 c0_U113:B 0 9.72738e-16
C189 c0_U10:Y 0 8.1474e-16
C190 c0_U68:B 0 2.78846e-16
C191 c0_U59:B 0 5.89356e-16
C192 c0_n10:9 0 1.66333e-15
C193 c0_n10:11 0 6.46572e-16
R138 c0_U115:A c0_U113:B 49.9471
R139 c0_U115:A c0_n10:9 35.0774
R140 c0_U113:B c0_n10:9 45.7227
R141 c0_U10:Y c0_n10:9 10
R142 c0_U68:B c0_n10:11 23.8667
R143 c0_U59:B c0_n10:9 12.3755
R144 c0_U59:B c0_n10:11 8.78939
R145 c0_n10:9 c0_n10:11 386.733
C194 iDFF_16_q_reg:Q 0 8.02749e-16
C195 c0_U170:A 0 3.19001e-16
C196 c0_U121:A 0 5.64383e-16
C197 c0_U58:A 0 4.66551e-16
C198 IN_N61:6 0 1.3495e-15
R146 iDFF_16_q_reg:Q IN_N61:6 74.7709
R147 iDFF_16_q_reg:Q c0_U58:A 35.0711
R148 c0_U58:A IN_N61:6 65.7583
R149 c0_U121:A IN_N61:6 7.73333
R150 c0_U121:A c0_U170:A 1.06667
C199 DFF_12_q_reg:D 0 6.139e-16
C200 c0_U67:Y 0 3.29517e-16
R151 c0_U67:Y DFF_12_q_reg:D 29.5333
C201 DFF_15_q_reg:D 0 6.57144e-16
C202 c0_U60:Y 0 3.35314e-16
R152 c0_U60:Y DFF_15_q_reg:D 28.7333
C203 oDFF_12_q_reg:D 0 5.38963e-16
C204 DFF_12_q_reg:Q 0 3.29546e-16
R153 DFF_12_q_reg:Q oDFF_12_q_reg:D 27.5333
C205 c0_U61:Y 0 1.60602e-16
C206 c0_U60:B 0 1.37487e-16
R154 c0_U61:Y c0_U60:B 0.866667
C207 c0_U68:Y 0 1.75503e-16
C208 c0_U67:B 0 1.25254e-15
R155 c0_U68:Y c0_U67:B 30.1333
C209 DFF_15_q_reg:CLK 0 5.07776e-16
C210 iDFF_12_q_reg:CLK 0 7.90749e-16
C211 oDFF_12_q_reg:CLK 0 4.26576e-16
C212 oDFF_14_q_reg:CLK 0 1.96819e-16
C213 oDFF_16_q_reg:CLK 0 8.60661e-16
C214 DFF_12_q_reg:CLK 0 9.19521e-16
C215 DFF_16_q_reg:CLK 0 3.67087e-16
C216 DFF_14_q_reg:CLK 0 4.29302e-16
C217 oDFF_11_q_reg:CLK 0 7.31603e-16
C218 oDFF_3_q_reg:CLK 0 4.77416e-16
C219 DFF_3_q_reg:CLK 0 3.28087e-16
C220 clk__L2_I2:Y 0 3.20368e-16
C221 DFF_7_q_reg:CLK 0 1.33354e-15
C222 oDFF_6_q_reg:CLK 0 2.23438e-16
C223 iDFF_7_q_reg:CLK 0 3.72759e-16
C224 oDFF_2_q_reg:CLK 0 2.62409e-16
C225 DFF_4_q_reg:CLK 0 1.20305e-16
C226 DFF_1_q_reg:CLK 0 3.42883e-16
C227 oDFF_1_q_reg:CLK 0 3.87377e-16
C228 oDFF_4_q_reg:CLK 0 4.76376e-16
C229 iDFF_4_q_reg:CLK 0 3.62752e-16
C230 DFF_5_q_reg:CLK 0 5.53606e-16
C231 DFF_2_q_reg:CLK 0 3.76326e-16
C232 iDFF_8_q_reg:CLK 0 5.38072e-16
C233 iDFF_14_q_reg:CLK 0 3.24364e-16
C234 DFF_15_q_reg:CLK 0 1.27826e-16
C235 oDFF_15_q_reg:CLK 0 7.55972e-16
C236 oDFF_15_q_reg:CLK 0 3.00984e-16
C237 oDFF_11_q_reg:CLK 0 3.69985e-16
C238 DFF_11_q_reg:CLK 0 7.38238e-16
C239 oDFF_3_q_reg:CLK 0 3.71212e-16
C240 iDFF_2_q_reg:CLK 0 1.52117e-16
C241 oDFF_7_q_reg:CLK 0 4.74871e-16
C242 oDFF_7_q_reg:CLK 0 3.06151e-16
C243 DFF_8_q_reg:CLK 0 6.53649e-16
C244 oDFF_8_q_reg:CLK 0 6.75942e-16
C245 iDFF_4_q_reg:CLK 0 2.56177e-16
C246 clk__L2_N2:52 0 1.18108e-15
C247 clk__L2_N2:75 0 8.79326e-16
C248 clk__L2_N2:81 0 2.28323e-15
C249 clk__L2_N2:89 0 2.20541e-15
R156 DFF_15_q_reg:CLK iDFF_12_q_reg:CLK 56.5773
R157 oDFF_12_q_reg:CLK DFF_15_q_reg:CLK 706.663
R158 DFF_15_q_reg:CLK DFF_12_q_reg:CLK 868.607
R159 oDFF_11_q_reg:CLK DFF_15_q_reg:CLK 212.396
R160 oDFF_3_q_reg:CLK DFF_15_q_reg:CLK 2925.38
R161 DFF_15_q_reg:CLK DFF_3_q_reg:CLK 4051.44
R162 oDFF_15_q_reg:CLK DFF_15_q_reg:CLK 81.5198
R163 DFF_15_q_reg:CLK DFF_11_q_reg:CLK 151.847
R164 DFF_15_q_reg:CLK clk__L2_N2:89 1406.75
R165 oDFF_12_q_reg:CLK iDFF_12_q_reg:CLK 178.176
R166 DFF_12_q_reg:CLK iDFF_12_q_reg:CLK 219.008
R167 oDFF_11_q_reg:CLK iDFF_12_q_reg:CLK 277.35
R168 oDFF_3_q_reg:CLK iDFF_12_q_reg:CLK 3820.01
R169 DFF_3_q_reg:CLK iDFF_12_q_reg:CLK 5290.45
R170 oDFF_15_q_reg:CLK iDFF_12_q_reg:CLK 20.5541
R171 DFF_11_q_reg:CLK iDFF_12_q_reg:CLK 198.284
R172 iDFF_12_q_reg:CLK clk__L2_N2:89 1836.96
R173 oDFF_12_q_reg:CLK DFF_12_q_reg:CLK 36.0303
R174 oDFF_12_q_reg:CLK oDFF_11_q_reg:CLK 3464.17
R175 oDFF_12_q_reg:CLK oDFF_3_q_reg:CLK 47712.8
R176 oDFF_12_q_reg:CLK DFF_3_q_reg:CLK 66078.9
R177 oDFF_15_q_reg:CLK oDFF_12_q_reg:CLK 118.258
R178 oDFF_12_q_reg:CLK DFF_11_q_reg:CLK 2476.61
R179 oDFF_12_q_reg:CLK clk__L2_N2:89 22944.1
R180 oDFF_16_q_reg:CLK oDFF_14_q_reg:CLK 35.9887
R181 oDFF_14_q_reg:CLK DFF_16_q_reg:CLK 99.3754
R182 oDFF_14_q_reg:CLK DFF_14_q_reg:CLK 118.526
R183 oDFF_16_q_reg:CLK DFF_16_q_reg:CLK 113.868
R184 oDFF_16_q_reg:CLK DFF_14_q_reg:CLK 135.811
R185 oDFF_16_q_reg:CLK DFF_12_q_reg:CLK 42.6
R186 oDFF_11_q_reg:CLK DFF_12_q_reg:CLK 4258.04
R187 oDFF_3_q_reg:CLK DFF_12_q_reg:CLK 58646.9
R188 DFF_12_q_reg:CLK DFF_3_q_reg:CLK 81222
R189 oDFF_15_q_reg:CLK DFF_12_q_reg:CLK 145.359
R190 DFF_12_q_reg:CLK DFF_11_q_reg:CLK 3044.17
R191 DFF_12_q_reg:CLK clk__L2_N2:89 28202.1
R192 DFF_16_q_reg:CLK DFF_14_q_reg:CLK 36.989
R193 oDFF_11_q_reg:CLK oDFF_3_q_reg:CLK 190.154
R194 oDFF_11_q_reg:CLK DFF_3_q_reg:CLK 263.35
R195 oDFF_15_q_reg:CLK oDFF_11_q_reg:CLK 399.622
R196 oDFF_11_q_reg:CLK DFF_11_q_reg:CLK 19.0526
R197 oDFF_11_q_reg:CLK clk__L2_N2:89 91.441
R198 oDFF_3_q_reg:CLK DFF_3_q_reg:CLK 126.936
R199 oDFF_15_q_reg:CLK oDFF_3_q_reg:CLK 5504.09
R200 oDFF_3_q_reg:CLK DFF_11_q_reg:CLK 262.415
R201 oDFF_3_q_reg:CLK clk__L2_N2:89 44.0752
R202 oDFF_15_q_reg:CLK DFF_3_q_reg:CLK 7622.78
R203 DFF_11_q_reg:CLK DFF_3_q_reg:CLK 363.427
R204 DFF_3_q_reg:CLK clk__L2_N2:89 36.3504
R205 DFF_7_q_reg:CLK clk__L2_I2:Y 145.362
R206 clk__L2_I2:Y clk__L2_N2:75 18.1298
R207 DFF_7_q_reg:CLK clk__L2_N2:75 42.3972
R208 DFF_7_q_reg:CLK iDFF_7_q_reg:CLK 86.3008
R209 oDFF_7_q_reg:CLK DFF_7_q_reg:CLK 117.765
R210 DFF_7_q_reg:CLK clk__L2_N2:89 29.2602
R211 oDFF_6_q_reg:CLK clk__L2_N2:75 28.8667
R212 oDFF_7_q_reg:CLK iDFF_7_q_reg:CLK 19.939
R213 iDFF_7_q_reg:CLK clk__L2_N2:89 38.3559
R214 oDFF_2_q_reg:CLK DFF_2_q_reg:CLK 237.998
R215 oDFF_2_q_reg:CLK iDFF_8_q_reg:CLK 215.124
R216 oDFF_2_q_reg:CLK DFF_8_q_reg:CLK 915.465
R217 oDFF_8_q_reg:CLK oDFF_2_q_reg:CLK 1336.3
R218 oDFF_2_q_reg:CLK clk__L2_N2:81 5122.47
R219 oDFF_2_q_reg:CLK clk__L2_N2:89 30.1733
R220 DFF_4_q_reg:CLK clk__L2_N2:81 12.8
R221 oDFF_1_q_reg:CLK DFF_1_q_reg:CLK 139.153
R222 oDFF_4_q_reg:CLK DFF_1_q_reg:CLK 136.477
R223 DFF_1_q_reg:CLK iDFF_4_q_reg:CLK 113.608
R224 DFF_5_q_reg:CLK DFF_1_q_reg:CLK 182.36
R225 DFF_1_q_reg:CLK clk__L2_N2:81 85.1489
R226 oDFF_4_q_reg:CLK oDFF_1_q_reg:CLK 40.6569
R227 oDFF_1_q_reg:CLK iDFF_4_q_reg:CLK 182.432
R228 oDFF_1_q_reg:CLK DFF_5_q_reg:CLK 292.835
R229 oDFF_1_q_reg:CLK clk__L2_N2:81 136.732
R230 oDFF_4_q_reg:CLK iDFF_4_q_reg:CLK 178.924
R231 oDFF_4_q_reg:CLK DFF_5_q_reg:CLK 287.203
R232 oDFF_4_q_reg:CLK clk__L2_N2:81 134.103
R233 DFF_5_q_reg:CLK iDFF_4_q_reg:CLK 204.334
R234 iDFF_4_q_reg:CLK clk__L2_N2:81 95.4089
R235 DFF_5_q_reg:CLK clk__L2_N2:81 35.6991
R236 DFF_2_q_reg:CLK iDFF_8_q_reg:CLK 52.0717
R237 DFF_8_q_reg:CLK DFF_2_q_reg:CLK 159.339
R238 oDFF_8_q_reg:CLK DFF_2_q_reg:CLK 232.586
R239 DFF_2_q_reg:CLK clk__L2_N2:81 891.579
R240 DFF_2_q_reg:CLK clk__L2_N2:89 57.8468
R241 DFF_8_q_reg:CLK iDFF_8_q_reg:CLK 200.295
R242 oDFF_8_q_reg:CLK iDFF_8_q_reg:CLK 292.369
R243 iDFF_8_q_reg:CLK clk__L2_N2:81 1120.75
R244 iDFF_8_q_reg:CLK clk__L2_N2:89 52.2872
R245 iDFF_14_q_reg:CLK clk__L2_N2:52 24.6
R246 DFF_15_q_reg:CLK clk__L2_N2:52 6.73333
R247 oDFF_15_q_reg:CLK DFF_11_q_reg:CLK 285.699
R248 oDFF_15_q_reg:CLK clk__L2_N2:89 2646.8
R249 oDFF_15_q_reg:CLK iDFF_16_q_reg:CLK 0.8
R250 oDFF_11_q_reg:CLK iDFF_11_q_reg:CLK 1.06667
R251 DFF_11_q_reg:CLK clk__L2_N2:89 126.19
R252 oDFF_3_q_reg:CLK iDFF_15_q_reg:CLK 1.06667
R253 iDFF_2_q_reg:CLK clk__L2_N2:75 13.1333
R254 oDFF_7_q_reg:CLK clk__L2_N2:89 52.3398
R255 oDFF_7_q_reg:CLK iDFF_3_q_reg:CLK 0.8
R256 oDFF_8_q_reg:CLK DFF_8_q_reg:CLK 19.5169
R257 DFF_8_q_reg:CLK clk__L2_N2:81 74.8149
R258 DFF_8_q_reg:CLK clk__L2_N2:89 222.509
R259 oDFF_8_q_reg:CLK clk__L2_N2:81 51.7125
R260 oDFF_8_q_reg:CLK clk__L2_N2:89 324.794
R261 iDFF_4_q_reg:CLK iDFF_1_q_reg:CLK 0.666667
R262 clk__L2_N2:81 clk__L2_N2:89 1245.05
C250 iDFF_5_q_reg:D 0 1.66398e-16
C251 N17 0 3.3063e-15
C252 N17:4 0 2.25136e-15
R263 iDFF_5_q_reg:D N17:4 14
R264 N17 N17:4 14.7167
C253 DFF_1_q_reg:D 0 1.97385e-15
C254 c0_U93:Y 0 2.3534e-16
R265 c0_U93:Y DFF_1_q_reg:D 32.3333
C255 DFF_5_q_reg:D 0 7.19973e-16
C256 c0_U83:Y 0 1.07496e-16
R266 c0_U83:Y DFF_5_q_reg:D 15.4
C257 oDFF_5_q_reg:D 0 1.01614e-15
C258 DFF_5_q_reg:Q 0 5.71834e-16
R267 DFF_5_q_reg:Q oDFF_5_q_reg:D 29.4667
C259 iDFF_33_q_reg:D 0 1.84928e-16
C260 N129 0 3.40929e-15
C261 N129:4 0 9.15052e-16
R268 iDFF_33_q_reg:D N129:4 10.3333
R269 N129 N129:4 43.9833
C262 N132 0 3.86421e-15
C263 iDFF_36_q_reg:D 0 1.31512e-16
R270 N132 iDFF_36_q_reg:D 24.5167
C264 N137 0 2.23452e-15
C265 iDFF_41_q_reg:D 0 1.42993e-16
C266 N137:2 0 1.90113e-15
R271 N137 N137:2 24.5833
R272 iDFF_41_q_reg:D N137:2 12.7333
C267 c0_U122:Y 0 1.86114e-16
C268 c0_U118:A 0 4.50566e-16
C269 c0_n98:3 0 2.82379e-15
R273 c0_U122:Y c0_n98:3 29.6
R274 c0_U118:A c0_n98:3 8.4
C270 iDFF_40_q_reg:Q 0 2.26256e-16
R275 iDFF_40_q_reg:Q c0_U110:A 0.8
C271 c0_U110:Y 0 3.4986e-16
R276 c0_U110:Y c0_U109:A 1.06667
C272 c0_U123:Y 0 6.72723e-16
C273 c0_U122:A 0 5.72785e-16
R277 c0_U123:Y c0_U122:A 15.7333
C274 c0_U131:Y 0 8.65109e-16
C275 c0_U130:A 0 2.14323e-16
R278 c0_U131:Y c0_U130:A 16
C276 c0_U177:Y 0 5.04341e-16
C277 c0_U173:A 0 8.79891e-16
R279 c0_U177:Y c0_U173:A 28.0667
C278 c0_U181:Y 0 6.75309e-16
C279 c0_U177:A 0 1.83682e-15
R280 c0_U181:Y c0_U177:A 31.8
C280 iDFF_6_q_reg:D 0 1.19175e-16
C281 N21 0 4.98438e-16
C282 N21:3 0 1.11667e-15
C283 N21:4 0 3.29024e-15
R281 iDFF_6_q_reg:D N21:3 8.06667
R282 N21 N21:4 10.1167
R283 N21:3 N21:4 51.4
C284 iDFF_34_q_reg:D 0 1.62325e-16
C285 N130 0 1.92906e-15
C286 N130:4 0 4.74863e-15
C287 N130:6 0 2.01129e-15
R284 iDFF_34_q_reg:D N130:6 14
R285 N130 N130:4 11.7167
R286 N130:4 N130:6 29.6667
C288 iDFF_40_q_reg:D 0 1.2981e-16
C289 N136 0 1.71898e-16
C290 N136:3 0 5.62067e-16
C291 N136:4 0 3.50336e-15
R287 iDFF_40_q_reg:D N136:3 8.4
R288 N136 N136:4 7.38333
R289 N136:3 N136:4 48.4667
C292 c0_U95:Y 0 1.80806e-16
C293 c0_U90:B 0 4.58948e-16
C294 c0_U88:B 0 5.0213e-16
C295 c0_U94:B 0 2.63527e-16
C296 c0_U92:B 0 5.98476e-16
C297 c0_n74:5 0 5.55618e-16
C298 c0_n74:7 0 1.40906e-15
C299 c0_n74:10 0 2.65662e-15
C300 c0_n74:12 0 3.31372e-15
R290 c0_U95:Y c0_n74:12 32.8
R291 c0_U90:B c0_n74:12 24.4667
R292 c0_U88:B c0_n74:5 9.06667
R293 c0_U94:B c0_n74:7 14.6811
R294 c0_U94:B c0_n74:10 27.16
R295 c0_U92:B c0_n74:10 17.6
R296 c0_n74:5 c0_n74:7 18.6667
R297 c0_n74:7 c0_n74:10 15.6692
R298 c0_n74:10 c0_n74:12 19.8667
C301 c0_U84:B 0 1.00951e-15
C302 c0_U80:B 0 8.715e-17
C303 c0_U78:B 0 1.47611e-16
C304 c0_U82:B 0 7.73343e-17
C305 c0_U85:Y 0 3.26909e-16
C306 c0_n68:5 0 8.73861e-16
C307 c0_n68:6 0 9.58305e-16
C308 c0_n68:10 0 2.14293e-15
C309 c0_n68:11 0 1.24343e-15
R299 c0_U84:B c0_n68:10 58.4417
R300 c0_U84:B c0_n68:11 27.502
R301 c0_U80:B c0_n68:5 9.73333
R302 c0_U78:B c0_n68:10 13.4667
R303 c0_U82:B c0_n68:6 6.81294
R304 c0_U82:B c0_n68:11 547.76
R305 c0_U85:Y c0_n68:6 39.1333
R306 c0_n68:5 c0_n68:10 23.2
R307 c0_n68:6 c0_n68:11 28.5292
R308 c0_n68:10 c0_n68:11 15.7817
C310 c0_U158:B 0 3.42574e-16
C311 iDFF_6_q_reg:Q 0 1.19509e-15
C312 c0_U135:B 0 1.80747e-16
C313 iDFF_6_q_reg:Q 0 2.37599e-16
C314 c0_U81:A 0 6.97961e-16
C315 IN_N21:6 0 1.75883e-15
C316 IN_N21:8 0 6.14688e-16
R309 c0_U158:B IN_N21:8 8.33333
R310 iDFF_6_q_reg:Q c0_U81:A 47.0957
R311 iDFF_6_q_reg:Q IN_N21:6 67.7
R312 c0_U135:B IN_N21:6 17.4667
R313 iDFF_6_q_reg:Q IN_N21:8 20.8
R314 c0_U81:A IN_N21:6 18.0533
C317 c0_U112:A 0 6.00041e-16
C318 c0_U34:C 0 1.73902e-16
C319 c0_U84:A 0 9.10937e-16
C320 c0_U173:Y 0 3.10752e-16
C321 c0_U7:A 0 1.09009e-16
C322 c0_U94:A 0 1.32295e-15
C323 c0_U173:Y 0 6.21235e-16
C324 c0_n30:10 0 1.6891e-15
C325 c0_n30:15 0 2.98385e-15
R315 c0_U112:A c0_n30:10 25.7648
R316 c0_U112:A c0_n30:15 61.1141
R317 c0_U34:C c0_n30:10 27.7333
R318 c0_U173:Y c0_U84:A 30.7333
R319 c0_U173:Y c0_n30:15 7.73333
R320 c0_U7:A c0_n30:10 7.4
R321 c0_U94:A c0_n30:15 23.7333
R322 c0_n30:10 c0_n30:15 159.151
C326 c0_U167:Y 0 2.40804e-16
C327 c0_U165:A 0 5.79769e-16
R323 c0_U167:Y c0_U165:A 15
C328 c0_U82:A 0 1.53954e-16
C329 c0_U114:C 0 2.06565e-16
C330 c0_U92:A 0 6.18331e-17
C331 c0_U132:A 0 5.65938e-17
C332 c0_U8:A 0 1.23067e-16
C333 c0_U133:Y 0 6.57551e-16
C334 c0_n62:8 0 1.53872e-15
C335 c0_n62:11 0 2.28944e-15
C336 c0_n62:15 0 1.01272e-15
C337 c0_n62:16 0 7.42713e-16
R324 c0_U82:A c0_n62:11 165.333
R325 c0_U82:A c0_n62:15 15.0303
R326 c0_U114:C c0_n62:16 13.8667
R327 c0_U92:A c0_n62:11 6.4
R328 c0_U132:A c0_n62:8 6.4
R329 c0_U8:A c0_n62:16 13.7333
R330 c0_U133:Y c0_n62:11 35.6667
R331 c0_n62:8 c0_n62:15 28.6667
R332 c0_n62:8 c0_n62:16 14.3333
R333 c0_n62:11 c0_n62:15 13.7778
C338 c0_U95:A 0 6.62094e-16
C339 c0_U85:A 0 6.59686e-16
C340 c0_U1:Y 0 7.45964e-16
R334 c0_U1:Y c0_U85:A 34.2937
R335 c0_U1:Y c0_U95:A 75.2747
R336 c0_U85:A c0_U95:A 69.6988
C341 c0_U132:Y 0 5.86074e-16
C342 c0_U111:A 0 9.16574e-16
C343 c0_U6:A 0 5.23607e-16
R337 c0_U132:Y c0_U6:A 51.1104
R338 c0_U132:Y c0_U111:A 17.4557
R339 c0_U6:A c0_U111:A 62.6353
C344 c0_U81:B 0 1.9786e-16
R340 c0_U82:Y c0_U81:B 0.533333
C345 c0_U112:Y 0 8.13015e-16
C346 c0_U111:C 0 1.3563e-15
R341 c0_U112:Y c0_U111:C 18.5333
C347 c0_U141:Y 0 3.85075e-16
C348 c0_U137:A 0 1.53167e-16
R342 c0_U141:Y c0_U137:A 1.4
C349 c0_U145:Y 0 5.95745e-16
C350 c0_U141:A 0 4.60895e-16
R343 c0_U145:Y c0_U141:A 15.4333
C351 c0_U165:B 0 2.81433e-16
C352 c0_U166:Y 0 1.36683e-16
C353 c0_n140:2 0 1.57449e-15
C354 c0_n140:5 0 1.75418e-15
R344 c0_U165:B c0_n140:5 21.7333
R345 c0_U166:Y c0_n140:2 7.06667
R346 c0_n140:2 c0_n140:5 14.2
C355 c0_U176:Y 0 5.51205e-16
C356 c0_U174:A 0 8.71246e-16
C357 c0_n146:4 0 2.8316e-15
R347 c0_U176:Y c0_n146:4 50.6667
R348 c0_U174:A c0_n146:4 15.7333
C358 iDFF_10_q_reg:Q 0 1.14934e-15
C359 c0_U167:B 0 3.05172e-16
C360 c0_U135:A 0 1.24044e-15
C361 c0_U71:A 0 4.6429e-16
C362 IN_N37:8 0 1.72565e-15
R349 iDFF_10_q_reg:Q c0_U71:A 31.1333
R350 iDFF_10_q_reg:Q c0_U167:B 0.8
R351 c0_U167:B IN_N37:8 11.6667
R352 c0_U135:A IN_N37:8 25.3333
C363 c0_U61:A 0 1.6374e-16
C364 c0_U59:A 0 7.22045e-17
C365 c0_U63:A 0 7.16832e-16
C366 c0_U66:Y 0 3.15492e-16
C367 c0_U65:A 0 6.48646e-16
C368 c0_n54:8 0 8.01082e-16
C369 c0_n54:12 0 3.20513e-15
R353 c0_U61:A c0_U59:A 421.067
R354 c0_U61:A c0_n54:8 21.0533
R355 c0_U59:A c0_n54:8 7.11261
R356 c0_U65:A c0_U63:A 16.5333
R357 c0_U63:A c0_n54:8 26.2
R358 c0_U66:Y c0_n54:12 26.2667
R359 c0_U65:A c0_n54:12 12.7333
C370 c0_U70:A 0 8.38792e-16
C371 c0_U74:A 0 1.00255e-15
C372 c0_U68:A 0 1.53047e-16
C373 c0_U75:Y 0 4.17895e-16
C374 c0_U72:A 0 3.02577e-16
C375 c0_n59:6 0 2.16813e-15
R360 c0_U70:A c0_n59:6 10.7333
R361 c0_U74:A c0_U72:A 3.2
R362 c0_U74:A c0_n59:6 30.4
R363 c0_U68:A c0_n59:6 8.73333
R364 c0_U75:Y c0_U72:A 29.0667
C376 iDFF_10_q_reg:D 0 2.34642e-15
C377 N37 0 6.2975e-17
C378 N37:2 0 4.01648e-15
C379 N37:3 0 5.42975e-16
R365 iDFF_10_q_reg:D N37:3 16.4
R366 N37 N37:2 18.45
R367 N37:2 N37:3 28.9333
C380 iDFF_38_q_reg:D 0 3.5254e-16
C381 N134 0 1.19993e-16
C382 N134:3 0 3.02215e-15
C383 N134:6 0 2.19357e-15
R368 iDFF_38_q_reg:D N134:6 48.4667
R369 N134 N134:3 13.85
R370 N134:3 N134:6 21.6667
C384 iDFF_41_q_reg:Q 0 3.23281e-16
C385 c0_U124:B 0 4.4662e-16
C386 c0_U110:B 0 5.99536e-16
C387 c0_U145:B 0 5.40252e-16
C388 c0_U159:B 0 1.42575e-15
C389 c0_U103:B 0 7.57043e-16
C390 c0_U185:B 0 4.09796e-16
C391 c0_U131:B 0 7.74419e-16
C392 c0_U172:A 0 4.85925e-16
C393 IN_N137:16 0 1.61405e-15
C394 IN_N137:19 0 1.08743e-15
C395 IN_N137:20 0 1.03242e-15
R371 iDFF_41_q_reg:Q c0_U124:B 49.5333
R372 iDFF_41_q_reg:Q IN_N137:19 56.227
R373 c0_U124:B IN_N137:19 18.575
R374 c0_U110:B IN_N137:20 15.8
R375 c0_U145:B IN_N137:20 16
R376 c0_U159:B c0_U103:B 78.3314
R377 c0_U185:B c0_U159:B 41.1741
R378 c0_U172:A c0_U159:B 41.2056
R379 c0_U159:B IN_N137:16 21.7747
R380 c0_U159:B IN_N137:20 53.9418
R381 c0_U185:B c0_U103:B 2617.96
R382 c0_U172:A c0_U103:B 82.3831
R383 c0_U103:B IN_N137:16 1384.5
R384 c0_U103:B IN_N137:20 107.847
R385 c0_U185:B c0_U172:A 1377.16
R386 c0_U185:B IN_N137:16 12.9256
R387 c0_U185:B IN_N137:20 1802.82
R388 c0_U131:B IN_N137:19 15.4667
R389 c0_U172:A IN_N137:16 728.303
R390 c0_U172:A IN_N137:20 23.5965
R391 IN_N137:16 IN_N137:19 9.6
R392 IN_N137:16 IN_N137:20 953.415
C396 c0_U116:Y 0 6.96728e-16
C397 c0_U114:A 0 9.13276e-17
C398 c0_U24:B 0 3.3538e-16
C399 c0_U43:A 0 4.80199e-16
C400 c0_n21:7 0 3.86408e-15
R393 c0_U116:Y c0_n21:7 18
R394 c0_U114:A c0_n21:7 15.8
R395 c0_U43:A c0_U24:B 19.1857
R396 c0_U24:B c0_n21:7 53.72
R397 c0_U43:A c0_n21:7 45.1084
C401 c0_U52:A 0 6.70104e-16
C402 c0_U114:B 0 7.08734e-17
C403 c0_U33:A 0 1.98223e-16
C404 c0_U115:Y 0 4.61732e-16
C405 c0_n27:5 0 1.81045e-15
R398 c0_U52:A c0_U33:A 19.19
R399 c0_U52:A c0_n27:5 61.5402
R400 c0_U115:Y c0_U114:B 160.32
R401 c0_U114:B c0_n27:5 7.70769
R402 c0_U33:A c0_n27:5 54.4936
R403 c0_U115:Y c0_n27:5 25.05
C406 c0_U52:B 0 5.68514e-17
C407 c0_U43:B 0 8.72572e-17
C408 c0_U53:Y 0 5.13843e-16
C409 c0_U34:B 0 1.10079e-16
C410 c0_n29:4 0 5.59677e-16
C411 c0_n29:6 0 3.36043e-16
C412 c0_n29:9 0 5.31878e-16
R404 c0_U52:B c0_n29:4 6.4
R405 c0_U43:B c0_n29:9 12.8
R406 c0_U53:Y c0_n29:9 19.8667
R407 c0_U34:B c0_n29:6 7.06667
R408 c0_n29:4 c0_n29:6 17.4
R409 c0_n29:4 c0_n29:9 8.53333
C413 c0_U85:C 0 2.24801e-16
C414 c0_U86:Y 0 2.3068e-16
C415 c0_U56:A 0 1.72535e-16
C416 c0_U66:B 0 7.13211e-17
C417 c0_n51:8 0 1.35435e-15
C418 c0_n51:9 0 1.30113e-15
R410 c0_U85:C c0_n51:9 21.5333
R411 c0_U86:Y c0_U56:A 17.7836
R412 c0_U86:Y c0_n51:8 64.8361
R413 c0_U56:A c0_n51:8 46.4498
R414 c0_U66:B c0_n51:8 6.4
R415 c0_n51:8 c0_n51:9 6
C419 c0_U95:C 0 9.50025e-16
C420 c0_U56:B 0 3.71725e-16
C421 c0_U75:A 0 2.54145e-16
C422 c0_U96:Y 0 3.21399e-16
C423 c0_n52:8 0 1.65462e-15
R416 c0_U95:C c0_n52:8 19.1333
R417 c0_U96:Y c0_U56:B 55.5312
R418 c0_U56:B c0_n52:8 28.6911
R419 c0_U75:A c0_n52:8 27.8667
R420 c0_U96:Y c0_n52:8 34.0884
C424 c0_U85:B 0 1.66714e-16
C425 c0_U111:Y 0 6.24664e-16
C426 c0_U95:B 0 1.08082e-16
C427 c0_U76:B 0 1.32902e-16
C428 c0_n65:5 0 1.83498e-15
C429 c0_n65:6 0 4.67644e-16
R421 c0_U111:Y c0_U85:B 53.6
R422 c0_U85:B c0_n65:5 26.8
R423 c0_U111:Y c0_n65:5 31.825
R424 c0_U95:B c0_n65:5 8.73333
R425 c0_U76:B c0_n65:6 8.06667
R426 c0_n65:5 c0_n65:6 34.5333
C430 c0_U101:B 0 4.34553e-16
C431 c0_U164:B 0 8.07292e-17
C432 c0_U165:Y 0 3.31769e-16
C433 c0_n83:5 0 1.90728e-15
C434 c0_n83:7 0 1.75431e-15
R427 c0_U101:B c0_n83:5 22.0667
R428 c0_U164:B c0_n83:5 6.4
R429 c0_U165:Y c0_n83:7 14.7333
R430 c0_n83:5 c0_n83:7 46.0267
C435 c0_U168:B 0 1.2465e-15
C436 c0_U169:Y 0 1.39338e-16
C437 c0_U108:B 0 1.51372e-15
C438 c0_n91:5 0 2.33013e-15
R431 c0_U168:B c0_U108:B 31.8
R432 c0_U169:Y c0_n91:5 6.73333
R433 c0_U108:B c0_n91:5 58.24
C439 c0_U72:B 0 2.64369e-17
C440 c0_U34:A 0 5.58563e-16
C441 c0_U8:Y 0 1.65966e-15
C442 c0_U63:B 0 5.08216e-16
C443 c0_n8:5 0 5.81773e-16
C444 c0_n8:6 0 1.68293e-15
R434 c0_U72:B c0_n8:5 58.7298
R435 c0_U72:B c0_n8:6 35.8032
R436 c0_U34:A c0_n8:5 8.4
R437 c0_U8:Y c0_n8:6 11.7333
R438 c0_U63:B c0_n8:6 8.8
R439 c0_n8:5 c0_n8:6 69.7417
C445 oDFF_20_q_reg:CLK 0 3.30649e-16
C446 DFF_24_q_reg:CLK 0 3.32536e-16
C447 DFF_20_q_reg:CLK 0 3.09343e-16
C448 iDFF_24_q_reg:CLK 0 2.27607e-16
C449 iDFF_23_q_reg:CLK 0 1.8518e-16
C450 oDFF_24_q_reg:CLK 0 7.3535e-16
C451 oDFF_5_q_reg:CLK 0 8.31548e-17
C452 iDFF_41_q_reg:CLK 0 8.69508e-16
C453 iDFF_5_q_reg:CLK 0 1.42276e-16
C454 iDFF_35_q_reg:CLK 0 5.3959e-16
C455 iDFF_36_q_reg:CLK 0 7.10961e-16
C456 iDFF_37_q_reg:CLK 0 3.85117e-16
C457 iDFF_20_q_reg:CLK 0 2.06077e-16
C458 iDFF_33_q_reg:CLK 0 8.32124e-17
C459 DFF_6_q_reg:CLK 0 2.46622e-16
C460 iDFF_6_q_reg:CLK 0 8.20284e-16
C461 iDFF_40_q_reg:CLK 0 6.75487e-16
C462 iDFF_13_q_reg:CLK 0 1.85366e-15
C463 iDFF_10_q_reg:CLK 0 2.35088e-16
C464 iDFF_38_q_reg:CLK 0 1.57676e-15
C465 iDFF_34_q_reg:CLK 0 5.98061e-16
C466 iDFF_31_q_reg:CLK 0 9.5695e-16
C467 DFF_31_q_reg:CLK 0 1.68539e-16
C468 iDFF_32_q_reg:CLK 0 7.29872e-16
C469 oDFF_32_q_reg:CLK 0 6.89464e-16
C470 oDFF_13_q_reg:CLK 0 3.70717e-16
C471 DFF_13_q_reg:CLK 0 8.17298e-16
C472 oDFF_9_q_reg:CLK 0 1.94068e-16
C473 oDFF_10_q_reg:CLK 0 5.9772e-16
C474 DFF_28_q_reg:CLK 0 4.87312e-16
C475 iDFF_9_q_reg:CLK 0 5.75225e-16
C476 DFF_32_q_reg:CLK 0 1.76017e-16
C477 DFF_10_q_reg:CLK 0 1.79453e-16
C478 DFF_9_q_reg:CLK 0 4.51868e-16
C479 iDFF_23_q_reg:CLK 0 2.71344e-16
C480 iDFF_6_q_reg:CLK 0 4.53033e-16
C481 clk__L2_I1:Y 0 3.45904e-16
C482 DFF_31_q_reg:CLK 0 1.75191e-16
C483 oDFF_9_q_reg:CLK 0 1.24701e-16
C484 oDFF_10_q_reg:CLK 0 2.92358e-16
C485 oDFF_28_q_reg:CLK 0 4.2847e-16
C486 clk__L2_N1:61 0 1.16057e-15
C487 clk__L2_N1:64 0 2.08712e-15
C488 clk__L2_N1:70 0 1.73753e-15
C489 clk__L2_N1:74 0 9.90603e-16
C490 clk__L2_N1:76 0 1.1687e-15
C491 clk__L2_N1:79 0 5.68804e-16
C492 clk__L2_N1:84 0 5.83034e-16
C493 clk__L2_N1:85 0 9.90575e-16
R440 oDFF_20_q_reg:CLK clk__L2_N1:61 28.2
R441 DFF_24_q_reg:CLK clk__L2_N1:61 13.0667
R442 DFF_24_q_reg:CLK DFF_20_q_reg:CLK 510.298
R443 DFF_24_q_reg:CLK iDFF_41_q_reg:CLK 39.69
R444 DFF_24_q_reg:CLK iDFF_37_q_reg:CLK 170.162
R445 DFF_24_q_reg:CLK iDFF_20_q_reg:CLK 671.445
R446 DFF_24_q_reg:CLK clk__L2_N1:70 83.9306
R447 DFF_20_q_reg:CLK iDFF_41_q_reg:CLK 520.111
R448 DFF_20_q_reg:CLK iDFF_37_q_reg:CLK 316.659
R449 DFF_20_q_reg:CLK iDFF_20_q_reg:CLK 175.59
R450 DFF_20_q_reg:CLK clk__L2_N1:70 21.9488
R451 oDFF_24_q_reg:CLK iDFF_24_q_reg:CLK 93.8583
R452 iDFF_24_q_reg:CLK iDFF_23_q_reg:CLK 68.7817
R453 iDFF_23_q_reg:CLK clk__L2_N1:61 17.3333
R454 oDFF_24_q_reg:CLK iDFF_23_q_reg:CLK 16.6859
R455 oDFF_5_q_reg:CLK clk__L2_N1:64 12.8
R456 iDFF_41_q_reg:CLK iDFF_36_q_reg:CLK 37.7546
R457 iDFF_41_q_reg:CLK clk__L2_N1:64 51.9953
R458 iDFF_41_q_reg:CLK iDFF_37_q_reg:CLK 173.434
R459 iDFF_41_q_reg:CLK iDFF_20_q_reg:CLK 684.357
R460 iDFF_41_q_reg:CLK clk__L2_N1:70 85.5446
R461 iDFF_5_q_reg:CLK clk__L2_N1:64 32.2
R462 iDFF_36_q_reg:CLK iDFF_35_q_reg:CLK 27.4667
R463 iDFF_36_q_reg:CLK clk__L2_N1:64 60.4844
R464 iDFF_37_q_reg:CLK iDFF_20_q_reg:CLK 416.657
R465 iDFF_37_q_reg:CLK clk__L2_N1:70 52.0821
R466 iDFF_20_q_reg:CLK clk__L2_N1:70 16.7712
R467 iDFF_33_q_reg:CLK clk__L2_N1:70 12.8
R468 DFF_6_q_reg:CLK iDFF_6_q_reg:CLK 42.4
R469 iDFF_40_q_reg:CLK clk__L2_N1:84 21.3333
R470 iDFF_13_q_reg:CLK iDFF_10_q_reg:CLK 32
R471 iDFF_10_q_reg:CLK clk__L2_N1:76 12.8
R472 iDFF_38_q_reg:CLK clk__L2_N1:76 41
R473 iDFF_34_q_reg:CLK clk__L2_I1:Y 14.4667
R474 iDFF_34_q_reg:CLK clk__L2_N1:84 23.4667
R475 DFF_31_q_reg:CLK iDFF_31_q_reg:CLK 16.4667
R476 DFF_31_q_reg:CLK iDFF_32_q_reg:CLK 27.4667
R477 DFF_28_q_reg:CLK iDFF_32_q_reg:CLK 56.4152
R478 oDFF_28_q_reg:CLK iDFF_32_q_reg:CLK 76.9833
R479 iDFF_32_q_reg:CLK clk__L2_N1:74 56.7894
R480 oDFF_32_q_reg:CLK clk__L2_N1:74 13.8667
R481 oDFF_32_q_reg:CLK clk__L2_N1:85 22.1333
R482 oDFF_13_q_reg:CLK DFF_13_q_reg:CLK 72.6267
R483 oDFF_13_q_reg:CLK iDFF_9_q_reg:CLK 66.0242
R484 DFF_13_q_reg:CLK iDFF_9_q_reg:CLK 35.0853
R485 DFF_13_q_reg:CLK clk__L2_N1:79 28.2
R486 oDFF_9_q_reg:CLK clk__L2_N1:79 16.2667
R487 oDFF_10_q_reg:CLK oDFF_9_q_reg:CLK 14.8
R488 oDFF_28_q_reg:CLK DFF_28_q_reg:CLK 18.7456
R489 DFF_28_q_reg:CLK clk__L2_N1:74 80.7512
R490 DFF_32_q_reg:CLK clk__L2_N1:74 13.3333
R491 DFF_10_q_reg:CLK DFF_9_q_reg:CLK 291.973
R492 DFF_10_q_reg:CLK clk__L2_N1:85 22.6922
R493 DFF_9_q_reg:CLK clk__L2_N1:85 30.4139
R494 iDFF_40_q_reg:CLK iDFF_6_q_reg:CLK 1.33333
R495 iDFF_38_q_reg:CLK clk__L2_I1:Y 0.8
R496 oDFF_10_q_reg:CLK DFF_28_q_reg:CLK 0.8
R497 oDFF_28_q_reg:CLK clk__L2_N1:74 110.192
R498 clk__L2_N1:70 clk__L2_N1:84 16.2
R499 clk__L2_N1:76 clk__L2_N1:85 11
C494 clk__L2_I1:A 0 1.04939e-16
C495 clk__L2_I2:A 0 5.50588e-15
C496 clk__L1_I0:Y 0 1.48095e-16
C497 clk__L2_I0:A 0 1.25661e-16
C498 clk__L1_N0:6 0 1.55325e-15
C499 clk__L1_N0:7 0 5.13091e-15
R500 clk__L2_I1:A clk__L2_I2:A 205.333
R501 clk__L2_I1:A clk__L1_N0:7 16.2105
R502 clk__L2_I2:A clk__L1_N0:7 38.5
R503 clk__L1_I0:Y clk__L1_N0:6 13.0667
R504 clk__L2_I0:A clk__L1_N0:7 33.6
R505 clk__L1_N0:6 clk__L1_N0:7 34.4667
C500 c0_U49:B 0 4.93726e-16
C501 c0_U51:B 0 1.32636e-16
C502 c0_U45:B 0 2.48596e-16
C503 c0_U47:B 0 9.01412e-16
C504 c0_U52:Y 0 1.98395e-16
C505 c0_n41:7 0 2.22183e-15
C506 c0_n41:11 0 2.12651e-15
R506 c0_U51:B c0_U49:B 20.0267
R507 c0_U49:B c0_U47:B 1.62159
R508 c0_U51:B c0_U47:B 100.133
R509 c0_U45:B c0_n41:7 7.6
R510 c0_U47:B c0_n41:7 29.2667
R511 c0_U52:Y c0_n41:11 34.6
R512 c0_n41:7 c0_n41:11 16.8667
C507 c0_U142:Y 0 1.38879e-16
C508 c0_U122:B 0 1.19093e-15
C509 c0_U141:B 0 3.72232e-16
C510 c0_n103:5 0 1.70796e-15
C511 c0_n103:6 0 2.65226e-15
R513 c0_U142:Y c0_n103:6 35.7333
R514 c0_U122:B c0_n103:5 10.9333
R515 c0_U141:B c0_n103:5 21
R516 c0_U141:B c0_n103:6 14
R517 c0_n103:5 c0_n103:6 10.9375
C512 c0_U146:Y 0 1.32535e-16
C513 c0_U53:A 0 4.99067e-16
C514 c0_U1:A 0 2.25375e-16
C515 c0_n46:6 0 9.98099e-16
C516 c0_n46:7 0 1.06474e-15
R518 c0_U146:Y c0_n46:7 25.6
R519 c0_U53:A c0_n46:6 28.3333
R520 c0_U53:A c0_n46:7 6.73333
R521 c0_U1:A c0_n46:6 7.26667
C517 c0_U129:B 0 3.46024e-16
C518 c0_U137:B 0 9.54773e-16
C519 c0_U138:Y 0 3.78892e-16
C520 c0_n111:3 0 1.61345e-15
C521 c0_n111:4 0 1.72532e-15
R522 c0_U129:B c0_n111:3 7.06667
R523 c0_U137:B c0_n111:3 41.1253
R524 c0_U137:B c0_n111:4 16.5828
R525 c0_U138:Y c0_n111:4 35.0667
R526 c0_n111:3 c0_n111:4 38.7975
C522 clk 0 3.22701e-15
C523 clk__L1_I0:A 0 2.86533e-16
R527 clk clk__L1_I0:A 47.45
C524 N29 0 2.83509e-15
C525 iDFF_8_q_reg:D 0 1.51453e-16
R528 N29 iDFF_8_q_reg:D 27.2333
C526 N33 0 2.98085e-16
C527 iDFF_9_q_reg:D 0 3.92272e-16
C528 N33:2 0 4.0332e-15
R529 N33 N33:2 40.7167
R530 iDFF_9_q_reg:D N33:2 14.8667
C529 iDFF_9_q_reg:Q 0 1.1581e-16
C530 c0_U176:B 0 8.82145e-16
C531 c0_U167:A 0 6.92647e-16
C532 c0_U73:A 0 5.54773e-16
C533 IN_N33:5 0 8.74981e-16
C534 IN_N33:9 0 1.37255e-15
R531 iDFF_9_q_reg:Q IN_N33:5 8.4
R532 c0_U73:A IN_N33:5 22
R533 c0_U73:A IN_N33:9 10.4
R534 c0_U167:A IN_N33:9 34.2341
R535 c0_U167:A c0_U176:B 18.941
R536 c0_U176:B IN_N33:9 48.1417
C535 DFF_14_q_reg:D 0 3.61796e-16
C536 c0_U62:Y 0 7.91836e-16
R537 c0_U62:Y DFF_14_q_reg:D 28.7333
C537 DFF_16_q_reg:D 0 3.84331e-16
C538 c0_U58:Y 0 6.70526e-16
R538 c0_U58:Y DFF_16_q_reg:D 30.6
C539 oDFF_14_q_reg:D 0 4.20268e-16
C540 DFF_14_q_reg:Q 0 3.86878e-16
R539 DFF_14_q_reg:Q oDFF_14_q_reg:D 28.1333
C541 oDFF_16_q_reg:D 0 1.40325e-16
C542 DFF_16_q_reg:Q 0 6.46035e-16
R540 DFF_16_q_reg:Q oDFF_16_q_reg:D 15.6
C543 c0_U63:Y 0 5.00019e-16
C544 c0_U62:B 0 2.76847e-16
R541 c0_U63:Y c0_U62:B 15.1333
C545 N41 0 2.12054e-15
C546 iDFF_11_q_reg:D 0 1.91298e-16
C547 N41:2 0 1.85875e-15
R542 N41 N41:2 11.8333
R543 iDFF_11_q_reg:D N41:2 19.8
C548 N45 0 3.05373e-15
C549 iDFF_12_q_reg:D 0 1.75991e-16
R544 N45 iDFF_12_q_reg:D 27.2333
C550 N49 0 2.16901e-15
C551 iDFF_13_q_reg:D 0 2.02309e-16
C552 N49:2 0 1.49189e-15
C553 N49:4 0 2.74233e-15
R545 N49 N49:4 12.1
R546 iDFF_13_q_reg:D N49:2 17.8667
R547 N49:2 N49:4 14.7333
C554 N53 0 3.70963e-15
C555 iDFF_14_q_reg:D 0 3.57185e-16
R548 N53 iDFF_14_q_reg:D 37.1883
C556 N57 0 2.11932e-15
C557 iDFF_15_q_reg:D 0 1.7796e-16
C558 N57:2 0 1.86281e-15
R549 N57 N57:2 11.8333
R550 iDFF_15_q_reg:D N57:2 19.8
C559 N61 0 3.81694e-15
C560 iDFF_16_q_reg:D 0 1.51453e-16
R551 N61 iDFF_16_q_reg:D 30.4333
C561 Qout_N726 0 1.25611e-15
C562 oDFF_3_q_reg:Q 0 2.05765e-15
R552 oDFF_3_q_reg:Q Qout_N726 26.4333
C563 Qout_N734 0 1.25611e-15
C564 oDFF_11_q_reg:Q 0 2.05765e-15
R553 oDFF_11_q_reg:Q Qout_N734 26.4333
C565 Qout_N735 0 1.25611e-15
C566 oDFF_12_q_reg:Q 0 2.04184e-15
R554 oDFF_12_q_reg:Q Qout_N735 26.4333
C567 Qout_N738 0 1.25546e-15
C568 oDFF_15_q_reg:Q 0 1.96596e-15
R555 oDFF_15_q_reg:Q Qout_N738 26.1667
C569 N77 0 4.40636e-15
C570 iDFF_20_q_reg:D 0 1.47026e-16
R556 N77 iDFF_20_q_reg:D 28.1833
C571 N133 0 2.22919e-16
C572 iDFF_37_q_reg:D 0 2.66828e-16
C573 N133:3 0 5.67297e-15
R557 N133 N133:3 6.93333
R558 iDFF_37_q_reg:D N133:3 38
C574 Qout_N724 0 1.57277e-15
C575 oDFF_1_q_reg:Q 0 1.15454e-16
C576 Qout_N724:3 0 1.99207e-15
R559 oDFF_1_q_reg:Q Qout_N724:3 13.0667
R560 Qout_N724 Qout_N724:3 7.38333
C577 Qout_N727 0 2.59069e-15
C578 oDFF_4_q_reg:Q 0 9.12481e-17
R561 oDFF_4_q_reg:Q Qout_N727 20.1833
C579 Qout_N733 0 2.8018e-17
C580 oDFF_10_q_reg:Q 0 9.43659e-16
C581 Qout_N733:2 0 2.98706e-15
R562 oDFF_10_q_reg:Q Qout_N733:2 24.0667
R563 Qout_N733 Qout_N733:2 16.1167
C582 Qout_N736 0 7.15138e-17
C583 oDFF_13_q_reg:Q 0 1.11178e-15
C584 Qout_N736:2 0 2.72951e-15
R564 oDFF_13_q_reg:Q Qout_N736:2 12.2667
R565 Qout_N736 Qout_N736:2 11.7833
C585 Qout_N737 0 5.96796e-17
C586 oDFF_14_q_reg:Q 0 3.26975e-15
R566 oDFF_14_q_reg:Q Qout_N737 23.5167
C587 Qout_N755 0 5.96796e-17
C588 oDFF_32_q_reg:Q 0 1.14683e-15
C589 Qout_N755:2 0 3.01829e-15
C590 Qout_N755:3 0 8.47252e-16
R567 oDFF_32_q_reg:Q Qout_N755:3 10.7333
R568 Qout_N755 Qout_N755:2 16.1167
R569 Qout_N755:2 Qout_N755:3 32.2667
C591 iDFF_1_q_reg:Q 0 4.35656e-16
C592 c0_U175:B 0 2.0928e-16
C593 c0_U154:A 0 2.18757e-16
C594 c0_U93:A 0 2.00242e-15
R570 iDFF_1_q_reg:Q c0_U93:A 58.7333
R571 iDFF_1_q_reg:Q c0_U175:B 17.4802
R572 c0_U93:A c0_U154:A 17.6667
R573 c0_U93:A c0_U175:B 46.9867
C595 iDFF_13_q_reg:Q 0 4.28085e-16
C596 c0_U176:A 0 5.87944e-16
R574 iDFF_13_q_reg:Q c0_U13:A 0.8
R575 iDFF_13_q_reg:Q c0_U176:A 15
C597 iDFF_14_q_reg:Q 0 9.06433e-16
C598 c0_U171:B 0 4.39086e-16
C599 c0_U136:A 0 2.84894e-15
C600 c0_U62:A 0 3.84973e-16
R576 iDFF_14_q_reg:Q c0_U171:B 20.3671
R577 iDFF_14_q_reg:Q c0_U62:A 15.8
R578 iDFF_14_q_reg:Q c0_U136:A 49.0083
R579 c0_U136:A c0_U171:B 31.7892
C601 iDFF_33_q_reg:Q 0 5.36748e-16
C602 c0_U185:A 0 1.00936e-16
R580 iDFF_33_q_reg:Q c0_U185:A 14.4667
C603 c0_U145:A 0 4.83021e-16
R581 iDFF_34_q_reg:Q c0_U145:A 1.6
C604 iDFF_35_q_reg:Q 0 7.19825e-16
C605 c0_U131:A 0 6.46292e-16
R582 iDFF_35_q_reg:Q c0_U131:A 29.6
C606 c0_U124:Y 0 1.75497e-15
C607 c0_U123:A 0 1.51815e-16
R583 c0_U124:Y c0_U123:A 18.7333
C608 iDFF_36_q_reg:Q 0 1.54701e-16
R584 iDFF_36_q_reg:Q c0_U124:A 0.533333
C609 iDFF_38_q_reg:Q 0 1.53332e-16
C610 c0_U172:B 0 8.52973e-16
R585 iDFF_38_q_reg:Q c0_U172:B 15.4
C611 DFF_9_q_reg:D 0 2.67559e-16
C612 c0_U73:Y 0 1.46949e-15
R586 c0_U73:Y DFF_9_q_reg:D 30.6
C613 DFF_10_q_reg:D 0 1.71578e-16
C614 c0_U71:Y 0 7.32798e-16
R587 c0_U71:Y DFF_10_q_reg:D 27.7333
C615 c0_U65:Y 0 7.44349e-16
C616 c0_U64:B 0 2.0021e-16
R588 c0_U65:Y c0_U64:B 15.4333
C617 c0_U72:Y 0 1.25465e-15
C618 c0_U71:B 0 2.22554e-16
R589 c0_U72:Y c0_U71:B 17.3333
C619 c0_U74:Y 0 5.63691e-16
C620 c0_U73:B 0 1.892e-16
R590 c0_U74:Y c0_U73:B 15.0667
C621 DFF_13_q_reg:D 0 5.04595e-16
C622 c0_U64:Y 0 9.0904e-16
R591 c0_U64:Y DFF_13_q_reg:D 29.8
C623 oDFF_1_q_reg:D 0 5.69828e-16
C624 DFF_1_q_reg:Q 0 2.25443e-16
R592 DFF_1_q_reg:Q oDFF_1_q_reg:D 15.0667
C625 oDFF_3_q_reg:D 0 4.47029e-16
C626 DFF_3_q_reg:Q 0 7.71557e-16
R593 DFF_3_q_reg:Q oDFF_3_q_reg:D 29.2
C627 oDFF_6_q_reg:D 0 6.51947e-16
C628 DFF_6_q_reg:Q 0 2.16208e-16
R594 DFF_6_q_reg:Q oDFF_6_q_reg:D 27.7333
C629 oDFF_7_q_reg:D 0 8.24646e-16
C630 DFF_7_q_reg:Q 0 5.86699e-16
R595 DFF_7_q_reg:Q oDFF_7_q_reg:D 29.4667
C631 oDFF_8_q_reg:D 0 5.74126e-16
C632 DFF_8_q_reg:Q 0 3.56966e-16
R596 DFF_8_q_reg:Q oDFF_8_q_reg:D 28.6667
C633 oDFF_9_q_reg:D 0 7.22288e-16
C634 DFF_9_q_reg:Q 0 6.29317e-16
R597 DFF_9_q_reg:Q oDFF_9_q_reg:D 28.6667
C635 oDFF_10_q_reg:D 0 2.00837e-16
C636 DFF_10_q_reg:Q 0 1.2857e-16
C637 Q_N733:4 0 1.12462e-15
R598 DFF_10_q_reg:Q Q_N733:4 19.7333
R599 oDFF_10_q_reg:D Q_N733:4 10
C638 oDFF_13_q_reg:D 0 6.61864e-16
C639 DFF_13_q_reg:Q 0 3.93443e-16
R600 DFF_13_q_reg:Q oDFF_13_q_reg:D 28.6667
C640 oDFF_15_q_reg:D 0 7.33853e-16
C641 DFF_15_q_reg:Q 0 5.85231e-16
R601 DFF_15_q_reg:Q oDFF_15_q_reg:D 29.4667
C642 c0_U33:B 0 6.74289e-16
C643 c0_U24:A 0 6.37915e-16
C644 c0_U2:Y 0 4.15155e-16
R602 c0_U2:Y c0_U24:A 54.2428
R603 c0_U2:Y c0_U33:B 18.1954
R604 c0_U24:A c0_U33:B 45.9979
C645 c0_U75:B 0 3.18636e-16
C646 c0_U66:A 0 1.23863e-15
C647 c0_U4:Y 0 6.7843e-16
R605 c0_U4:Y c0_U66:A 57.0375
R606 c0_U4:Y c0_U75:B 41.9586
R607 c0_U66:A c0_U75:B 43.4571
C648 c0_U52:C 0 1.02585e-15
C649 c0_U43:C 0 2.2374e-16
C650 c0_U6:Y 0 6.31071e-16
R608 c0_U6:Y c0_U52:C 2.13333
R609 c0_U43:C c0_U52:C 27.2
C651 c0_U132:B 0 1.30121e-16
C652 c0_U74:B 0 8.78546e-16
C653 c0_U65:B 0 2.51777e-16
C654 c0_U7:Y 0 1.71332e-15
C655 c0_n7:6 0 1.58203e-15
R610 c0_U7:Y c0_n7:6 8.4
R611 c0_U7:Y c0_U65:B 18.4
R612 c0_U65:B c0_U74:B 3.2
R613 c0_U132:B c0_n7:6 22.4
C656 c0_U34:Y 0 7.478e-16
C657 c0_U2:A 0 6.44729e-16
R614 c0_U34:Y c0_U2:A 29.1333
C658 c0_U59:Y 0 8.00116e-16
C659 c0_U58:B 0 1.77505e-16
R615 c0_U59:Y c0_U58:B 15.1667
C660 c0_U152:Y 0 2.31965e-16
C661 c0_U151:B 0 3.3305e-16
C662 c0_U102:B 0 3.36233e-16
C663 c0_n85:4 0 3.30215e-15
R616 c0_U152:Y c0_n85:4 19.5333
R617 c0_U102:B c0_U151:B 1.06667
R618 c0_U151:B c0_n85:4 41.9067
C664 c0_U108:Y 0 7.40931e-16
C665 c0_U104:A 0 4.78477e-16
R619 c0_U108:Y c0_U104:A 3.8
C666 c0_U109:Y 0 3.18362e-15
C667 c0_U108:A 0 3.95345e-16
R620 c0_U109:Y c0_U108:A 23.2
C668 c0_U156:Y 0 3.79595e-16
C669 c0_U155:B 0 4.15877e-16
C670 c0_U109:B 0 4.13249e-16
C671 c0_n93:4 0 3.428e-15
R621 c0_U156:Y c0_n93:4 7.53333
R622 c0_U109:B c0_n93:4 30.5333
R623 c0_U109:B c0_U155:B 1.6
C672 c0_U117:Y 0 2.17347e-15
C673 c0_U111:B 0 3.1303e-16
R624 c0_U117:Y c0_U111:B 32.6
C674 c0_U114:Y 0 2.48569e-16
C675 c0_U113:C 0 9.42851e-16
R625 c0_U114:Y c0_U113:C 17
C676 c0_U182:Y 0 1.24268e-16
C677 c0_U181:B 0 1.68244e-16
C678 c0_U123:B 0 6.36005e-16
C679 c0_n105:3 0 2.71509e-15
R626 c0_U182:Y c0_n105:3 29.3333
R627 c0_U123:B c0_n105:3 8.33333
R628 c0_U181:B c0_n105:3 9.06667
C680 c0_U130:Y 0 7.11277e-16
C681 c0_U129:A 0 1.85173e-16
C682 c0_n110:3 0 1.63051e-15
C683 c0_n110:4 0 2.23634e-15
R629 c0_U130:Y c0_n110:4 8.73333
R630 c0_U129:A c0_n110:3 8.06667
R631 c0_n110:3 c0_n110:4 35.6667
C684 c0_U178:Y 0 1.28526e-16
C685 c0_U177:B 0 5.7898e-16
C686 c0_U130:B 0 1.33292e-15
C687 c0_n113:4 0 2.48948e-15
R632 c0_U178:Y c0_n113:4 25.6
R633 c0_U130:B c0_n113:4 31.0672
R634 c0_U130:B c0_U177:B 25.3385
R635 c0_U177:B c0_n113:4 24.4708
C688 c0_U172:Y 0 9.01041e-16
C689 c0_U168:A 0 1.87842e-16
R636 c0_U172:Y c0_U168:A 15.4333
C690 c0_U185:Y 0 8.54719e-16
C691 c0_U181:A 0 4.51853e-16
R637 c0_U185:Y c0_U181:A 28.8
C692 iDFF_39_q_reg:D 0 2.67473e-16
C693 N135 0 2.17408e-15
C694 N135:4 0 5.24161e-15
R638 iDFF_39_q_reg:D N135:4 26.9333
R639 N135 N135:4 24.7833
C695 N93 0 3.02992e-15
C696 iDFF_24_q_reg:D 0 1.2446e-16
C697 N93:2 0 9.31354e-16
R640 N93 N93:2 31.25
R641 iDFF_24_q_reg:D N93:2 9.73333
C698 Qout_N743 0 3.00171e-15
C699 oDFF_20_q_reg:Q 0 9.78161e-17
R642 oDFF_20_q_reg:Q Qout_N743 20.1833
C700 Qout_N746 0 2.59113e-15
C701 oDFF_23_q_reg:Q 0 9.40157e-17
R643 oDFF_23_q_reg:Q Qout_N746 20.1833
C702 Qout_N747 0 2.59069e-15
C703 oDFF_24_q_reg:Q 0 9.12481e-17
R644 oDFF_24_q_reg:Q Qout_N747 20.1833
C704 iDFF_24_q_reg:Q 0 2.36117e-16
C705 c0_U183:A 0 2.40228e-16
C706 c0_U107:A 0 1.50923e-16
C707 c0_U35:A 0 3.94234e-16
C708 IN_N93:4 0 1.59923e-15
R645 iDFF_24_q_reg:Q IN_N93:4 19.157
R646 iDFF_24_q_reg:Q c0_U183:A 86.6056
R647 c0_U35:A IN_N93:4 14.8
R648 c0_U107:A IN_N93:4 14.4667
R649 c0_U183:A IN_N93:4 21.2095
C709 c0_U103:A 0 5.53012e-16
R650 iDFF_39_q_reg:Q c0_U103:A 1.86667
C710 DFF_20_q_reg:D 0 5.67348e-16
C711 c0_U44:Y 0 2.5454e-16
R651 c0_U44:Y DFF_20_q_reg:D 15.6
C712 c0_U36:Y 0 2.88012e-16
C713 c0_U35:B 0 1.88317e-15
R652 c0_U36:Y c0_U35:B 19.9333
C714 c0_U38:Y 0 4.93509e-16
C715 c0_U37:B 0 1.96087e-15
R653 c0_U38:Y c0_U37:B 47
C716 c0_U45:Y 0 1.73919e-16
C717 c0_U44:B 0 1.56715e-15
R654 c0_U45:Y c0_U44:B 17.0667
C718 c0_U159:Y 0 9.2325e-16
C719 c0_U155:A 0 1.70519e-16
R655 c0_U159:Y c0_U155:A 16.5333
C720 c0_U179:Y 0 4.61216e-16
C721 c0_U178:B 0 8.09898e-16
R656 c0_U179:Y c0_U178:B 27.8
C722 c0_U184:Y 0 1.95713e-16
C723 c0_U182:A 0 4.06574e-16
C724 c0_n152:2 0 2.04118e-15
R657 c0_U184:Y c0_n152:2 28.3333
R658 c0_U182:A c0_n152:2 7.06667
C725 c0_U45:A 0 2.26058e-16
C726 c0_U104:Y 0 2.85816e-16
C727 c0_U57:B 0 3.38849e-16
C728 c0_U36:A 0 2.50457e-15
C729 c0_U11:A 0 2.00646e-16
C730 c0_U86:B 0 1.72047e-16
C731 c0_n32:9 0 9.97592e-16
C732 c0_n32:14 0 1.32364e-15
R659 c0_U57:B c0_U45:A 1800.17
R660 c0_U45:A c0_U36:A 29.0249
R661 c0_U45:A c0_n32:14 2587.75
R662 c0_U104:Y c0_n32:14 14.1333
R663 c0_U57:B c0_U36:A 34.6187
R664 c0_U57:B c0_n32:14 19.2219
R665 c0_U36:A c0_n32:14 49.7644
R666 c0_U11:A c0_n32:9 24.4923
R667 c0_U11:A c0_n32:14 22.7429
R668 c0_U86:B c0_n32:9 16.3333
R669 c0_n32:9 c0_n32:14 39.8
C733 c0_U19:Y 0 7.59866e-16
C734 c0_U18:B 0 1.90743e-16
R670 c0_U19:Y c0_U18:B 15.4667
C735 c0_U26:Y 0 1.71102e-15
C736 c0_U25:B 0 1.30197e-16
C737 c0_n22:2 0 1.02667e-15
R671 c0_U26:Y c0_n22:2 26.6667
R672 c0_U25:B c0_n22:2 8.06667
C738 c0_U57:Y 0 6.21883e-16
C739 c0_U53:B 0 1.61611e-16
R673 c0_U57:Y c0_U53:B 15.4
C740 c0_U53:C 0 4.27101e-16
R674 c0_U54:Y c0_U53:C 1.33333
C741 c0_U55:Y 0 1.58297e-16
C742 c0_U54:B 0 9.24061e-16
R675 c0_U55:Y c0_U54:B 15.1333
C743 c0_U76:Y 0 7.21874e-16
C744 c0_U4:A 0 2.07855e-16
C745 c0_n64:3 0 1.12901e-15
R676 c0_U76:Y c0_n64:3 15.6667
R677 c0_U4:A c0_n64:3 16
C746 c0_U98:Y 0 2.96933e-16
C747 c0_U97:B 0 5.66808e-16
R678 c0_U98:Y c0_U97:B 14.7333
C748 c0_U100:Y 0 5.24013e-16
C749 c0_U98:A 0 1.65539e-16
C750 c0_n80:3 0 1.51587e-15
C751 c0_n80:4 0 1.11391e-15
R679 c0_U100:Y c0_n80:4 8.73333
R680 c0_U98:A c0_n80:3 8.06667
R681 c0_n80:3 c0_n80:4 35.9333
C752 c0_U102:Y 0 6.21912e-16
C753 c0_U101:A 0 4.22532e-16
R682 c0_U102:Y c0_U101:A 27.5333
C754 c0_U103:Y 0 1.32696e-15
C755 c0_U102:A 0 2.41654e-16
R683 c0_U103:Y c0_U102:A 17.2
C756 c0_U105:Y 0 6.02633e-16
C757 c0_U104:B 0 4.22912e-16
R684 c0_U105:Y c0_U104:B 16
C758 c0_U106:Y 0 1.02696e-16
C759 c0_U105:B 0 1.83983e-15
C760 c0_n89:3 0 1.47853e-15
R685 c0_U106:Y c0_n89:3 10.7333
R686 c0_U105:B c0_n89:3 25.8
C761 c0_U139:Y 0 4.22104e-16
C762 c0_U138:B 0 2.20493e-16
R687 c0_U139:Y c0_U138:B 1.93333
C763 c0_U144:Y 0 1.33439e-16
C764 c0_U142:A 0 6.19663e-16
C765 c0_n122:2 0 1.18635e-15
R688 c0_U144:Y c0_n122:2 26.4
R689 c0_U142:A c0_n122:2 8.06667
C766 c0_U155:Y 0 7.06755e-16
C767 c0_U151:A 0 1.58169e-16
R690 c0_U155:Y c0_U151:A 15.7333
C768 c0_U168:Y 0 1.40303e-15
C769 c0_U164:A 0 3.68883e-16
R691 c0_U168:Y c0_U164:A 31.6
C770 iDFF_31_q_reg:D 0 1.45964e-15
C771 N121 0 7.06239e-17
C772 N121:2 0 3.73115e-15
R692 iDFF_31_q_reg:D N121:2 40
R693 N121 N121:2 17.1167
C773 iDFF_31_q_reg:Q 0 1.59241e-16
C774 c0_U143:B 0 3.6467e-16
C775 c0_U99:A 0 1.07867e-15
C776 c0_U18:A 0 1.32315e-15
R694 iDFF_31_q_reg:Q c0_U18:A 8.08333
R695 c0_U18:A c0_U143:B 26.6467
R696 c0_U18:A c0_U99:A 56.4357
R697 c0_U99:A c0_U143:B 93.8382
C777 DFF_28_q_reg:D 0 5.56543e-16
C778 c0_U25:Y 0 6.79442e-16
R698 c0_U25:Y DFF_28_q_reg:D 29.5333
C779 oDFF_28_q_reg:D 0 2.6448e-16
C780 DFF_28_q_reg:Q 0 4.284e-16
R699 DFF_28_q_reg:Q oDFF_28_q_reg:D 15.0667
C781 oDFF_31_q_reg:D 0 3.79934e-16
C782 DFF_31_q_reg:Q 0 5.6964e-16
R700 DFF_31_q_reg:Q oDFF_31_q_reg:D 28.4
C783 oDFF_32_q_reg:D 0 5.71347e-16
C784 DFF_32_q_reg:Q 0 1.80187e-16
R701 DFF_32_q_reg:Q oDFF_32_q_reg:D 26.9333
C785 c0_U17:Y 0 1.77589e-16
C786 c0_U16:B 0 1.41247e-16
R702 c0_U17:Y c0_U16:B 0.866667
C787 c0_U107:B 0 7.59727e-16
C788 c0_U179:A 0 2.58224e-16
C789 iDFF_20_q_reg:Q 0 6.75147e-16
C790 c0_U44:A 0 8.10295e-16
C791 IN_N77:4 0 2.05587e-15
R703 iDFF_20_q_reg:Q c0_U107:B 245.929
R704 c0_U107:B c0_U44:A 70.8986
R705 c0_U107:B IN_N77:4 12.1458
R706 c0_U179:A IN_N77:4 26.1333
R707 iDFF_20_q_reg:Q c0_U44:A 36.8363
R708 iDFF_20_q_reg:Q IN_N77:4 166.515
R709 c0_U44:A IN_N77:4 48.0042
C792 c0_U184:A 0 6.82797e-16
C793 iDFF_21_q_reg:Q 0 1.66888e-15
C794 c0_U150:B 0 4.54914e-16
C795 c0_U41:A 0 2.69499e-16
C796 IN_N81:8 0 2.01364e-15
C797 IN_N81:12 0 8.58785e-16
R710 c0_U184:A IN_N81:8 20.8
R711 iDFF_21_q_reg:Q IN_N81:8 13.2
R712 iDFF_21_q_reg:Q c0_U150:B 23.8053
R713 iDFF_21_q_reg:Q IN_N81:12 55.7938
R714 c0_U150:B IN_N81:12 29.2689
R715 c0_U41:A IN_N81:12 7.53333
C798 iDFF_18_q_reg:Q 0 6.16865e-16
C799 c0_U180:B 0 3.07512e-16
C800 c0_U163:B 0 3.76416e-16
C801 c0_U48:A 0 1.86991e-16
R716 iDFF_18_q_reg:Q c0_U163:B 1.33333
R717 iDFF_18_q_reg:Q c0_U180:B 47.4667
R718 iDFF_18_q_reg:Q c0_U48:A 23.7333
R719 c0_U48:A c0_U180:B 1.63678
C802 iDFF_22_q_reg:Q 0 5.46885e-16
C803 c0_U184:B 0 5.41673e-16
C804 c0_U163:A 0 4.09287e-16
R720 iDFF_22_q_reg:Q c0_U39:A 0.266667
R721 iDFF_22_q_reg:Q c0_U163:A 28.6
R722 c0_U163:A c0_U184:B 2.13333
C805 DFF_17_q_reg:D 0 7.04735e-16
C806 c0_U50:Y 0 7.56642e-16
R723 c0_U50:Y DFF_17_q_reg:D 30.3333
C807 DFF_22_q_reg:D 0 1.76876e-16
C808 c0_U39:Y 0 1.06272e-15
R724 c0_U39:Y DFF_22_q_reg:D 27.7333
C809 DFF_29_q_reg:D 0 2.91457e-16
C810 c0_U22:Y 0 1.32007e-16
C811 N752:2 0 1.19416e-15
R725 c0_U22:Y N752:2 6.73333
R726 DFF_29_q_reg:D N752:2 21.9333
C812 c0_U146:B 0 2.03528e-16
C813 c0_U32:B 0 2.49547e-16
C814 c0_U23:B 0 1.99209e-16
C815 c0_U3:Y 0 6.35824e-16
C816 c0_n3:4 0 2.38343e-15
R727 c0_U3:Y c0_n3:4 14.6667
R728 c0_U3:Y c0_U146:B 1.13333
R729 c0_U23:B c0_n3:4 14.2
R730 c0_U32:B c0_n3:4 19.6667
C817 c0_U180:A 0 3.7698e-16
C818 c0_U14:Y 0 2.42308e-16
R731 c0_U14:Y c0_U180:A 2.2
C819 c0_U23:Y 0 1.04753e-15
C820 c0_U22:B 0 2.50566e-16
R732 c0_U23:Y c0_U22:B 28
C821 c0_U47:Y 0 1.20086e-16
C822 c0_U46:B 0 2.44878e-15
C823 c0_n42:3 0 1.14283e-15
R733 c0_U47:Y c0_n42:3 7.06667
R734 c0_U46:B c0_n42:3 30.6
C824 c0_U51:Y 0 2.09201e-15
C825 c0_U50:B 0 3.86654e-16
R735 c0_U51:Y c0_U50:B 31.3333
C826 c0_U148:Y 0 4.11073e-16
C827 c0_U147:B 0 8.82483e-16
R736 c0_U148:Y c0_U147:B 28.3333
C828 c0_U150:Y 0 3.295e-16
C829 c0_U148:A 0 4.82786e-16
R737 c0_U150:Y c0_U148:A 27.8
C830 c0_U149:Y 0 3.64832e-16
C831 c0_U148:B 0 6.57979e-16
R738 c0_U149:Y c0_U148:B 27.2667
C832 c0_U161:Y 0 4.28754e-16
C833 c0_U160:B 0 8.55049e-16
R739 c0_U161:Y c0_U160:B 28.0667
C834 c0_U162:Y 0 1.10973e-16
C835 c0_U161:B 0 1.07413e-15
C836 c0_n137:4 0 1.22581e-15
R740 c0_U162:Y c0_n137:4 11.7333
R741 c0_U161:B c0_n137:4 35.5333
C837 c0_U97:Y 0 3.59239e-16
C838 c0_U57:A 0 2.8543e-16
C839 c0_U47:A 0 3.26374e-16
C840 c0_U5:A 0 1.76256e-17
C841 c0_U97:Y 0 1.40198e-16
C842 c0_U38:A 0 9.49467e-16
C843 c0_U96:B 0 9.63506e-17
C844 c0_n35:11 0 7.92734e-16
C845 c0_n35:14 0 3.91605e-16
C846 c0_n35:15 0 1.94849e-15
R742 c0_U97:Y c0_n35:14 14.8
R743 c0_U57:A c0_n35:15 14.8
R744 c0_U47:A c0_U38:A 27.2
R745 c0_U5:A c0_n35:11 25.2016
R746 c0_U5:A c0_n35:15 31.0078
R747 c0_U97:Y c0_U38:A 16.6
R748 c0_U96:B c0_n35:11 9.06667
R749 c0_n35:11 c0_n35:15 65.8917
R750 c0_n35:14 c0_n35:15 15
C847 c0_U106:A 0 8.83005e-16
C848 iDFF_32_q_reg:Q 0 9.6133e-17
C849 c0_U16:A 0 8.26926e-17
C850 c0_U143:A 0 4.35975e-16
C851 c0_U16:A 0 8.48729e-16
C852 IN_N125:6 0 2.39319e-15
R751 c0_U106:A IN_N125:6 13.3333
R752 iDFF_32_q_reg:Q c0_U16:A 11.15
R753 c0_U16:A IN_N125:6 6.4
R754 c0_U143:A IN_N125:6 25.3333
C853 c0_U55:A 0 1.62784e-16
C854 c0_U11:Y 0 9.59973e-16
C855 c0_U96:A 0 4.06613e-16
C856 c0_U17:B 0 4.90965e-16
C857 c0_U26:B 0 7.70818e-17
C858 c0_U11:Y 0 8.57496e-16
R755 c0_U55:A c0_U11:Y 29.6
R756 c0_U96:A c0_U11:Y 95.416
R757 c0_U17:B c0_U11:Y 137.823
R758 c0_U26:B c0_U11:Y 23.6401
R759 c0_U96:A c0_U17:B 21.4823
R760 c0_U96:A c0_U26:B 68.4006
R761 c0_U26:B c0_U17:B 98.8009
C859 c0_U23:A 0 7.14458e-16
C860 c0_U17:A 0 4.25746e-16
C861 c0_U21:A 0 1.76792e-15
C862 c0_U19:A 0 5.00562e-16
C863 c0_U24:Y 0 5.11144e-16
C864 c0_n17:9 0 2.55078e-15
C865 c0_n17:13 0 1.12062e-15
R762 c0_U23:A c0_U21:A 15.9333
R763 c0_U19:A c0_U17:A 121.953
R764 c0_U17:A c0_n17:13 14.6932
R765 c0_U21:A c0_n17:9 31.1333
R766 c0_U19:A c0_n17:9 6.73333
R767 c0_U19:A c0_n17:13 30.299
R768 c0_U24:Y c0_n17:13 23.4667
C866 iDFF_26_q_reg:Q 0 6.39584e-16
C867 c0_U162:B 0 5.09314e-16
C868 c0_U140:A 0 1.1095e-15
C869 c0_U29:A 0 4.73278e-16
R769 iDFF_26_q_reg:Q c0_U29:A 1.6
R770 iDFF_26_q_reg:Q c0_U140:A 66.6222
R771 iDFF_26_q_reg:Q c0_U162:B 19.4992
R772 c0_U140:A c0_U162:B 42.0772
C870 iDFF_30_q_reg:Q 0 5.04505e-16
C871 c0_U162:A 0 1.81092e-16
C872 c0_U15:A 0 3.72686e-16
C873 IN_N117:5 0 1.54396e-15
R773 iDFF_30_q_reg:Q IN_N117:5 24.8
R774 c0_U15:A IN_N117:5 8.66667
R775 c0_U162:A IN_N117:5 6.73333
C874 DFF_25_q_reg:D 0 1.55319e-16
C875 c0_U31:Y 0 2.29954e-16
C876 N748:2 0 1.25256e-15
R776 c0_U31:Y N748:2 7.06667
R777 DFF_25_q_reg:D N748:2 23.2
C877 DFF_30_q_reg:D 0 2.22883e-16
C878 c0_U20:Y 0 9.55559e-16
R778 c0_U20:Y DFF_30_q_reg:D 28.2667
C879 c0_U28:Y 0 1.12014e-15
C880 c0_U27:B 0 4.56361e-16
R779 c0_U28:Y c0_U27:B 18.0667
C881 c0_U38:B 0 2.5459e-16
C882 c0_U40:B 0 8.07009e-16
C883 c0_U42:B 0 5.79394e-17
C884 c0_U43:Y 0 9.98079e-16
C885 c0_U36:B 0 9.31505e-17
C886 c0_n33:10 0 1.75838e-15
C887 c0_n33:15 0 1.95837e-15
R780 c0_U40:B c0_U38:B 149.979
R781 c0_U38:B c0_n33:15 19.1208
R782 c0_U40:B c0_n33:15 21.236
R783 c0_U42:B c0_n33:10 6.4
R784 c0_U43:Y c0_n33:10 32.3333
R785 c0_U36:B c0_n33:15 15.9333
R786 c0_n33:10 c0_n33:15 27.8667
C888 c0_U40:A 0 6.32356e-16
C889 c0_U160:Y 0 4.30286e-16
C890 c0_U146:A 0 6.05227e-16
C891 c0_U49:A 0 2.11369e-16
C892 c0_U12:A 0 1.26872e-15
C893 c0_U56:C 0 2.3531e-16
C894 c0_n37:13 0 1.14921e-15
C895 c0_n37:16 0 1.19461e-15
R787 c0_U49:A c0_U40:A 19.4628
R788 c0_U40:A c0_n37:16 31.4243
R789 c0_U160:Y c0_U12:A 28.3333
R790 c0_U160:Y c0_n37:16 31.8667
R791 c0_U146:A c0_U12:A 17.2959
R792 c0_U146:A c0_n37:13 315.65
R793 c0_U49:A c0_n37:16 24.9317
R794 c0_U12:A c0_n37:13 27.8106
R795 c0_U56:C c0_n37:13 10.2667
C896 c0_U147:Y 0 3.3619e-16
C897 c0_U3:A 0 1.05571e-16
C898 c0_U42:A 0 7.6973e-17
C899 c0_U147:Y 0 6.02715e-16
C900 c0_U51:A 0 1.63144e-15
C901 c0_U76:C 0 7.80962e-17
C902 c0_U54:A 0 4.27415e-16
C903 c0_n39:11 0 9.70362e-16
C904 c0_n39:14 0 9.69047e-16
R796 c0_U147:Y c0_n39:11 24
R797 c0_U51:A c0_U3:A 19.1333
R798 c0_U42:A c0_n39:11 6.4
R799 c0_U147:Y c0_U51:A 14.8
R800 c0_U76:C c0_n39:14 8.73333
R801 c0_U54:A c0_n39:11 37.2
R802 c0_U54:A c0_n39:14 24.4667
C905 c0_U139:B 0 5.80686e-16
C906 c0_U106:B 0 3.53732e-16
C907 c0_U25:A 0 6.63779e-16
C908 iDFF_28_q_reg:Q 0 7.24368e-16
C909 IN_N109:6 0 3.43977e-15
R803 c0_U139:B IN_N109:6 28.2
R804 c0_U106:B IN_N109:6 7.66667
R805 iDFF_28_q_reg:Q c0_U25:A 60.1956
R806 c0_U25:A IN_N109:6 16.8773
R807 iDFF_28_q_reg:Q IN_N109:6 69.4564
C910 c0_U32:A 0 6.20186e-16
C911 c0_U30:A 0 4.58005e-16
C912 c0_U33:Y 0 4.22963e-16
C913 c0_U28:A 0 3.24658e-16
C914 c0_U26:A 0 2.34403e-16
C915 c0_n23:7 0 2.53707e-16
C916 c0_n23:9 0 3.26764e-15
R808 c0_U32:A c0_U30:A 38.4829
R809 c0_U32:A c0_U28:A 22.9463
R810 c0_U32:A c0_n23:9 68.1058
R811 c0_U30:A c0_U28:A 27.1868
R812 c0_U30:A c0_n23:9 118.103
R813 c0_U33:Y c0_n23:7 7.8
R814 c0_U28:A c0_n23:9 70.4214
R815 c0_U26:A c0_n23:9 8.2
R816 c0_n23:7 c0_n23:9 16.2667
C917 c0_U12:Y 0 1.08979e-16
C918 c0_U30:B 0 7.99508e-17
C919 c0_U76:A 0 1.55073e-16
C920 c0_U21:B 0 3.7126e-16
C921 c0_U12:Y 0 1.92047e-16
C922 c0_n12:7 0 9.34948e-16
C923 c0_n12:8 0 1.09882e-15
R817 c0_U12:Y c0_n12:8 29.6
R818 c0_U30:B c0_n12:7 13.7333
R819 c0_U76:A c0_n12:8 7
R820 c0_U21:B c0_U12:Y 0.8
R821 c0_U21:B c0_n12:7 9
C924 iDFF_27_q_reg:D 0 1.24833e-15
C925 N105 0 7.06239e-17
C926 N105:2 0 3.75666e-15
R822 iDFF_27_q_reg:D N105:2 39.6667
R823 N105 N105:2 17.45
C927 N109 0 7.06239e-17
C928 iDFF_28_q_reg:D 0 4.53628e-15
R824 N109 iDFF_28_q_reg:D 27.85
C929 Qout_N749 0 5.96796e-17
C930 oDFF_26_q_reg:Q 0 4.41592e-15
R825 oDFF_26_q_reg:Q Qout_N749 26.85
C931 DFF_27_q_reg:D 0 1.1313e-16
C932 c0_U27:Y 0 5.53408e-16
R826 c0_U27:Y DFF_27_q_reg:D 15.1333
C933 oDFF_26_q_reg:D 0 5.54293e-16
C934 DFF_26_q_reg:Q 0 3.16926e-16
R827 DFF_26_q_reg:Q oDFF_26_q_reg:D 28.7333
C935 oDFF_27_q_reg:D 0 2.26625e-16
C936 DFF_27_q_reg:Q 0 8.1916e-16
R828 DFF_27_q_reg:Q oDFF_27_q_reg:D 15.3333
C937 c0_U30:Y 0 7.30372e-16
R829 c0_U30:Y c0_U29:B 2.93333
C938 c0_U14:A 0 2.01826e-15
C939 c0_U50:A 0 1.88217e-16
C940 c0_U149:A 0 7.86857e-16
C941 iDFF_17_q_reg:Q 0 3.27253e-16
C942 IN_N65:6 0 1.76839e-15
R830 c0_U149:A c0_U14:A 28.2785
R831 c0_U14:A IN_N65:6 38.7237
R832 c0_U50:A IN_N65:6 13.8
R833 c0_U149:A IN_N65:6 23.7477
R834 iDFF_17_q_reg:Q IN_N65:6 17.3333
C943 c0_U150:A 0 1.15969e-15
C944 iDFF_25_q_reg:Q 0 8.76392e-16
C945 c0_U139:A 0 3.16052e-16
C946 c0_U31:A 0 2.75499e-16
C947 IN_N97:5 0 9.53432e-16
C948 IN_N97:7 0 2.19429e-15
C949 IN_N97:8 0 2.01622e-15
R835 c0_U150:A IN_N97:5 9.73333
R836 iDFF_25_q_reg:Q IN_N97:7 22.2
R837 c0_U139:A IN_N97:8 14.1333
R838 c0_U31:A IN_N97:7 14.3333
R839 c0_U31:A IN_N97:8 20.5333
R840 IN_N97:5 IN_N97:8 26.8667
C950 iDFF_21_q_reg:D 0 1.55793e-16
C951 N81 0 2.99376e-15
C952 N81:4 0 2.44284e-15
R841 iDFF_21_q_reg:D N81:4 6.73333
R842 N81 N81:4 29.9333
C953 iDFF_17_q_reg:CLK 0 1.73708e-16
C954 oDFF_17_q_reg:CLK 0 5.35202e-16
C955 DFF_18_q_reg:CLK 0 5.84838e-16
C956 iDFF_29_q_reg:CLK 0 2.98926e-16
C957 DFF_21_q_reg:CLK 0 9.176e-16
C958 iDFF_25_q_reg:CLK 0 1.47398e-16
C959 oDFF_30_q_reg:CLK 0 3.71839e-16
C960 oDFF_21_q_reg:CLK 0 7.01323e-16
C961 DFF_25_q_reg:CLK 0 6.59388e-16
C962 oDFF_26_q_reg:CLK 0 2.97146e-16
C963 DFF_26_q_reg:CLK 0 7.83708e-16
C964 iDFF_26_q_reg:CLK 0 1.33989e-16
C965 oDFF_25_q_reg:CLK 0 2.81842e-16
C966 oDFF_31_q_reg:CLK 0 2.50778e-16
C967 iDFF_28_q_reg:CLK 0 1.22639e-16
C968 DFF_27_q_reg:CLK 0 5.08516e-16
C969 oDFF_27_q_reg:CLK 0 3.5864e-16
C970 iDFF_27_q_reg:CLK 0 1.39779e-15
C971 oDFF_29_q_reg:CLK 0 2.68472e-16
C972 DFF_30_q_reg:CLK 0 2.45238e-16
C973 DFF_29_q_reg:CLK 0 1.45637e-16
C974 clk__L2_I0:Y 0 7.56796e-16
C975 iDFF_39_q_reg:CLK 0 1.31142e-15
C976 iDFF_21_q_reg:CLK 0 1.33027e-16
C977 DFF_17_q_reg:CLK 0 4.63314e-16
C978 iDFF_18_q_reg:CLK 0 1.19394e-16
C979 DFF_22_q_reg:CLK 0 2.61011e-16
C980 oDFF_22_q_reg:CLK 0 1.5073e-16
C981 DFF_19_q_reg:CLK 0 8.28432e-16
C982 iDFF_19_q_reg:CLK 0 1.37458e-15
C983 iDFF_22_q_reg:CLK 0 1.65319e-15
C984 oDFF_23_q_reg:CLK 0 8.43364e-16
C985 oDFF_17_q_reg:CLK 0 1.18208e-16
C986 iDFF_25_q_reg:CLK 0 3.04676e-16
C987 iDFF_25_q_reg:CLK 0 5.34918e-16
C988 iDFF_30_q_reg:CLK 0 6.52248e-16
C989 iDFF_26_q_reg:CLK 0 5.39856e-16
C990 iDFF_28_q_reg:CLK 0 4.2566e-16
C991 iDFF_21_q_reg:CLK 0 5.48987e-16
C992 iDFF_18_q_reg:CLK 0 5.3331e-16
C993 oDFF_19_q_reg:CLK 0 7.66012e-16
C994 DFF_19_q_reg:CLK 0 1.28702e-16
C995 DFF_23_q_reg:CLK 0 3.49195e-16
C996 clk__L2_N0:65 0 7.79643e-16
C997 clk__L2_N0:66 0 5.43608e-16
C998 clk__L2_N0:73 0 2.43257e-15
C999 clk__L2_N0:81 0 1.16247e-15
C1000 clk__L2_N0:84 0 1.0954e-15
C1001 clk__L2_N0:87 0 1.68415e-15
R843 iDFF_17_q_reg:CLK clk__L2_N0:84 22.1333
R844 oDFF_17_q_reg:CLK DFF_17_q_reg:CLK 61.1466
R845 oDFF_17_q_reg:CLK clk__L2_N0:84 47.7678
R846 oDFF_17_q_reg:CLK clk__L2_N0:87 66.2422
R847 oDFF_17_q_reg:CLK DFF_18_q_reg:CLK 14.8
R848 iDFF_29_q_reg:CLK iDFF_25_q_reg:CLK 18.3003
R849 iDFF_29_q_reg:CLK clk__L2_N0:84 30.551
R850 DFF_21_q_reg:CLK iDFF_25_q_reg:CLK 29.6
R851 oDFF_30_q_reg:CLK oDFF_21_q_reg:CLK 421.313
R852 oDFF_30_q_reg:CLK DFF_25_q_reg:CLK 136.412
R853 oDFF_30_q_reg:CLK oDFF_25_q_reg:CLK 1068.38
R854 oDFF_30_q_reg:CLK oDFF_29_q_reg:CLK 232.831
R855 oDFF_30_q_reg:CLK iDFF_30_q_reg:CLK 186.481
R856 oDFF_30_q_reg:CLK clk__L2_N0:73 58.2077
R857 oDFF_21_q_reg:CLK DFF_25_q_reg:CLK 839.424
R858 oDFF_25_q_reg:CLK oDFF_21_q_reg:CLK 6574.39
R859 oDFF_29_q_reg:CLK oDFF_21_q_reg:CLK 196.162
R860 oDFF_21_q_reg:CLK iDFF_30_q_reg:CLK 1147.53
R861 oDFF_21_q_reg:CLK clk__L2_N0:73 49.0405
R862 oDFF_25_q_reg:CLK DFF_25_q_reg:CLK 106.325
R863 oDFF_29_q_reg:CLK DFF_25_q_reg:CLK 463.892
R864 DFF_25_q_reg:CLK iDFF_30_q_reg:CLK 18.5586
R865 DFF_25_q_reg:CLK clk__L2_N0:73 115.973
R866 oDFF_26_q_reg:CLK DFF_26_q_reg:CLK 144.8
R867 oDFF_26_q_reg:CLK DFF_27_q_reg:CLK 40.596
R868 oDFF_27_q_reg:CLK oDFF_26_q_reg:CLK 100.058
R869 oDFF_26_q_reg:CLK iDFF_27_q_reg:CLK 199.927
R870 DFF_27_q_reg:CLK DFF_26_q_reg:CLK 150.37
R871 oDFF_27_q_reg:CLK DFF_26_q_reg:CLK 117.61
R872 DFF_26_q_reg:CLK iDFF_27_q_reg:CLK 44.0195
R873 DFF_26_q_reg:CLK clk__L2_N0:65 28.7333
R874 iDFF_26_q_reg:CLK clk__L2_N0:65 15.2
R875 oDFF_29_q_reg:CLK oDFF_25_q_reg:CLK 3633.22
R876 oDFF_25_q_reg:CLK iDFF_30_q_reg:CLK 76.2527
R877 oDFF_25_q_reg:CLK clk__L2_N0:73 908.304
R878 oDFF_31_q_reg:CLK clk__L2_N0:66 27.9333
R879 iDFF_28_q_reg:CLK clk__L2_N0:66 14.6667
R880 oDFF_27_q_reg:CLK DFF_27_q_reg:CLK 103.907
R881 DFF_27_q_reg:CLK iDFF_27_q_reg:CLK 207.617
R882 oDFF_27_q_reg:CLK iDFF_27_q_reg:CLK 162.385
R883 oDFF_29_q_reg:CLK iDFF_30_q_reg:CLK 634.161
R884 oDFF_29_q_reg:CLK clk__L2_N0:73 19.3127
R885 DFF_30_q_reg:CLK clk__L2_N0:73 27.8667
R886 DFF_29_q_reg:CLK clk__L2_I0:Y 511.467
R887 DFF_29_q_reg:CLK clk__L2_N0:73 13.9491
R888 clk__L2_I0:Y clk__L2_N0:73 31.9667
R889 iDFF_39_q_reg:CLK iDFF_21_q_reg:CLK 34.1333
R890 DFF_17_q_reg:CLK clk__L2_N0:84 42.5842
R891 DFF_17_q_reg:CLK clk__L2_N0:87 54.4122
R892 iDFF_18_q_reg:CLK clk__L2_N0:87 19.2
R893 DFF_22_q_reg:CLK iDFF_22_q_reg:CLK 64.354
R894 DFF_22_q_reg:CLK clk__L2_N0:81 67.7827
R895 DFF_22_q_reg:CLK clk__L2_N0:87 35.6057
R896 oDFF_22_q_reg:CLK clk__L2_N0:81 13.0667
R897 DFF_19_q_reg:CLK clk__L2_N0:81 15.4667
R898 oDFF_23_q_reg:CLK iDFF_19_q_reg:CLK 95.9076
R899 DFF_23_q_reg:CLK iDFF_19_q_reg:CLK 70.2835
R900 iDFF_22_q_reg:CLK iDFF_19_q_reg:CLK 29.0667
R901 iDFF_22_q_reg:CLK clk__L2_N0:81 86.1405
R902 iDFF_22_q_reg:CLK clk__L2_N0:87 45.2489
R903 oDFF_23_q_reg:CLK DFF_23_q_reg:CLK 16.6494
R904 iDFF_25_q_reg:CLK clk__L2_N0:84 38.5069
R905 oDFF_21_q_reg:CLK iDFF_25_q_reg:CLK 1.6
R906 iDFF_30_q_reg:CLK clk__L2_N0:73 158.54
R907 oDFF_25_q_reg:CLK iDFF_26_q_reg:CLK 1.6
R908 DFF_27_q_reg:CLK iDFF_28_q_reg:CLK 1.33333
R909 DFF_17_q_reg:CLK iDFF_21_q_reg:CLK 1.73333
R910 oDFF_18_q_reg:CLK iDFF_18_q_reg:CLK 1.6
R911 oDFF_19_q_reg:CLK DFF_19_q_reg:CLK 15.4
R912 clk__L2_N0:81 clk__L2_N0:87 47.6597
R913 clk__L2_N0:84 clk__L2_N0:87 46.1329
C1002 N65 0 3.15317e-15
C1003 iDFF_17_q_reg:D 0 1.87355e-16
R914 N65 iDFF_17_q_reg:D 27.7333
C1004 Qout_N744 0 1.25064e-15
C1005 oDFF_21_q_reg:Q 0 2.12074e-15
R915 oDFF_21_q_reg:Q Qout_N744 26.6667
C1006 Qout_N748 0 1.25064e-15
C1007 oDFF_25_q_reg:Q 0 2.11288e-15
R916 oDFF_25_q_reg:Q Qout_N748 26.6667
C1008 Qout_N752 0 1.25064e-15
C1009 oDFF_29_q_reg:Q 0 2.11288e-15
R917 oDFF_29_q_reg:Q Qout_N752 26.6667
C1010 Qout_N753 0 1.25064e-15
C1011 oDFF_30_q_reg:Q 0 2.11288e-15
R918 oDFF_30_q_reg:Q Qout_N753 26.6667
C1012 oDFF_25_q_reg:D 0 6.72098e-16
C1013 DFF_25_q_reg:Q 0 1.19894e-15
R919 DFF_25_q_reg:Q oDFF_25_q_reg:D 32.3333
C1014 N69 0 2.24133e-15
C1015 iDFF_18_q_reg:D 0 1.22108e-16
C1016 N69:4 0 1.82842e-15
R920 N69 N69:4 25.6667
R921 iDFF_18_q_reg:D N69:4 6.73333
C1017 Qout_N740 0 1.25064e-15
C1018 oDFF_17_q_reg:Q 0 2.11288e-15
R922 oDFF_17_q_reg:Q Qout_N740 26.6667
C1019 Qout_N741 0 1.25064e-15
C1020 oDFF_18_q_reg:Q 0 2.12376e-15
R923 oDFF_18_q_reg:Q Qout_N741 26.6667
C1021 oDFF_17_q_reg:D 0 2.39602e-16
C1022 DFF_17_q_reg:Q 0 9.83457e-16
R924 DFF_17_q_reg:Q oDFF_17_q_reg:D 27.7333
C1023 oDFF_18_q_reg:D 0 7.92351e-16
C1024 DFF_18_q_reg:Q 0 4.48006e-16
R925 DFF_18_q_reg:Q oDFF_18_q_reg:D 29.5333
C1025 oDFF_22_q_reg:D 0 9.56334e-16
C1026 DFF_22_q_reg:Q 0 3.09352e-16
R926 DFF_22_q_reg:Q oDFF_22_q_reg:D 29.5333
C1027 N73 0 2.94463e-15
C1028 iDFF_19_q_reg:D 0 1.14951e-16
C1029 N73:2 0 1.60827e-15
R927 N73 N73:2 42.05
R928 iDFF_19_q_reg:D N73:2 11.7333
C1030 N85 0 3.18707e-15
C1031 iDFF_22_q_reg:D 0 1.15358e-16
C1032 N85:2 0 1.81525e-15
R929 N85 N85:2 42.05
R930 iDFF_22_q_reg:D N85:2 11.7333
C1033 Qout_N745 0 3.4949e-16
C1034 oDFF_22_q_reg:Q 0 5.87566e-16
C1035 Qout_N745:3 0 3.29264e-15
R931 oDFF_22_q_reg:Q Qout_N745:3 43.6667
R932 Qout_N745 Qout_N745:3 7.46667
C1036 DFF_19_q_reg:D 0 6.52659e-16
C1037 c0_U46:Y 0 5.41766e-16
R933 c0_U46:Y DFF_19_q_reg:D 30.8667
C1038 oDFF_19_q_reg:D 0 8.8787e-16
C1039 DFF_19_q_reg:Q 0 2.93668e-16
R934 DFF_19_q_reg:Q oDFF_19_q_reg:D 29.2
C1040 oDFF_23_q_reg:D 0 6.07373e-16
C1041 DFF_23_q_reg:Q 0 3.74712e-16
R935 DFF_23_q_reg:Q oDFF_23_q_reg:D 28.6667
C1042 c0_U40:Y 0 5.16051e-16
C1043 c0_U39:B 0 5.0407e-16
C1044 c0_n36:2 0 3.21131e-15
R936 c0_U40:Y c0_n36:2 32.2667
R937 c0_U39:B c0_n36:2 33.6
C1045 N89 0 4.37721e-15
C1046 iDFF_23_q_reg:D 0 1.45243e-16
R938 N89 iDFF_23_q_reg:D 24.5167
C1047 N97 0 2.3313e-15
C1048 iDFF_25_q_reg:D 0 1.27863e-16
C1049 N97:4 0 1.7529e-15
R939 N97 N97:4 25.6667
R940 iDFF_25_q_reg:D N97:4 6.73333
C1050 N101 0 4.07552e-15
C1051 iDFF_26_q_reg:D 0 1.52501e-16
R941 N101 iDFF_26_q_reg:D 31.7333
C1052 N113 0 3.13827e-15
C1053 iDFF_29_q_reg:D 0 2.71963e-16
R942 N113 iDFF_29_q_reg:D 34.12
C1054 N117 0 3.18242e-15
C1055 iDFF_30_q_reg:D 0 1.67115e-16
R943 N117 iDFF_30_q_reg:D 28.8
C1056 N125 0 5.96796e-17
C1057 iDFF_32_q_reg:D 0 4.22487e-15
R944 N125 iDFF_32_q_reg:D 27.85
C1058 Qout_N732 0 5.96796e-17
C1059 oDFF_9_q_reg:Q 0 3.26358e-15
R945 oDFF_9_q_reg:Q Qout_N732 23.5167
C1060 Qout_N751 0 5.96796e-17
C1061 oDFF_28_q_reg:Q 0 3.26358e-15
R946 oDFF_28_q_reg:Q Qout_N751 23.5167
C1062 Qout_N742 0 2.85189e-15
C1063 oDFF_19_q_reg:Q 0 9.69547e-17
R947 oDFF_19_q_reg:Q Qout_N742 20.1833
C1064 Qout_N750 0 5.96796e-17
C1065 oDFF_27_q_reg:Q 0 3.26358e-15
R948 oDFF_27_q_reg:Q Qout_N750 23.5167
C1066 Qout_N754 0 7.06239e-17
C1067 oDFF_31_q_reg:Q 0 3.57872e-15
R949 oDFF_31_q_reg:Q Qout_N754 23.5167
C1068 iDFF_19_q_reg:Q 0 8.42874e-16
C1069 c0_U179:B 0 6.31272e-16
C1070 c0_U100:B 0 6.851e-16
R950 iDFF_19_q_reg:Q c0_U46:A 0.266667
R951 iDFF_19_q_reg:Q c0_U179:B 70.2673
R952 iDFF_19_q_reg:Q c0_U100:B 41.5783
R953 c0_U100:B c0_U179:B 21.3579
C1071 iDFF_23_q_reg:Q 0 1.06004e-15
C1072 c0_U183:B 0 4.15059e-16
C1073 c0_U100:A 0 2.15645e-16
C1074 c0_U37:A 0 4.50444e-16
R954 iDFF_23_q_reg:Q c0_U37:A 18.3764
R955 iDFF_23_q_reg:Q c0_U183:B 64.8917
R956 c0_U37:A c0_U183:B 44.4971
R957 c0_U100:A c0_U183:B 0.8
C1075 DFF_23_q_reg:D 0 2.12357e-16
C1076 c0_U37:Y 0 9.78992e-17
C1077 N746:2 0 8.77679e-16
R958 c0_U37:Y N746:2 8.73333
R959 DFF_23_q_reg:D N746:2 20
C1078 DFF_24_q_reg:D 0 3.0835e-16
C1079 c0_U35:Y 0 3.23889e-16
C1080 N747:2 0 1.01663e-15
R960 c0_U35:Y N747:2 24.9333
R961 DFF_24_q_reg:D N747:2 7.26667
C1081 oDFF_20_q_reg:D 0 4.52618e-16
C1082 DFF_20_q_reg:Q 0 1.13051e-16
C1083 Q_N743:3 0 9.16223e-16
R962 DFF_20_q_reg:Q Q_N743:3 10.7333
R963 oDFF_20_q_reg:D Q_N743:3 21.2667
C1084 iDFF_27_q_reg:Q 0 4.70732e-16
C1085 c0_U140:B 0 4.38466e-16
C1086 c0_U99:B 0 2.06142e-15
C1087 c0_U27:A 0 3.66212e-16
R964 iDFF_27_q_reg:Q c0_U99:B 23.8397
R965 iDFF_27_q_reg:Q c0_U27:A 39.85
R966 iDFF_27_q_reg:Q c0_U140:B 2503.16
R967 c0_U27:A c0_U99:B 78.4325
R968 c0_U27:A c0_U140:B 8235.41
R969 c0_U99:B c0_U140:B 28.6851
C1088 iDFF_29_q_reg:Q 0 2.25135e-16
C1089 c0_U149:B 0 2.52712e-16
C1090 c0_U144:A 0 3.95654e-16
C1091 c0_U22:A 0 3.30854e-16
C1092 IN_N113:4 0 1.25459e-15
C1093 IN_N113:5 0 1.36342e-15
R970 iDFF_29_q_reg:Q IN_N113:5 15.2
R971 c0_U22:A IN_N113:4 21.4
R972 c0_U144:A IN_N113:4 22.6667
R973 c0_U149:B IN_N113:5 13.0667
R974 IN_N113:4 IN_N113:5 12.7333
C1094 iDFF_37_q_reg:Q 0 6.39855e-16
C1095 c0_U159:A 0 4.03336e-16
R975 iDFF_37_q_reg:Q c0_U159:A 16.5333
C1096 DFF_18_q_reg:D 0 2.20925e-16
C1097 c0_U48:Y 0 1.11733e-15
R976 c0_U48:Y DFF_18_q_reg:D 29.0667
C1098 DFF_21_q_reg:D 0 2.81739e-16
C1099 c0_U41:Y 0 1.7531e-15
R977 c0_U41:Y DFF_21_q_reg:D 30.7333
C1100 DFF_26_q_reg:D 0 3.68101e-16
C1101 c0_U29:Y 0 4.01052e-16
R978 c0_U29:Y DFF_26_q_reg:D 15.3333
C1102 DFF_31_q_reg:D 0 5.03359e-16
C1103 c0_U18:Y 0 3.27617e-16
C1104 N754:3 0 1.66324e-15
R979 c0_U18:Y N754:3 20.4
R980 DFF_31_q_reg:D N754:3 25.5333
C1105 DFF_32_q_reg:D 0 9.29509e-16
C1106 c0_U16:Y 0 1.90654e-16
R981 c0_U16:Y DFF_32_q_reg:D 28
C1107 oDFF_21_q_reg:D 0 3.59989e-16
C1108 DFF_21_q_reg:Q 0 2.11232e-15
R982 DFF_21_q_reg:Q oDFF_21_q_reg:D 33.5333
C1109 oDFF_24_q_reg:D 0 1.24865e-15
C1110 DFF_24_q_reg:Q 0 1.39687e-15
R983 DFF_24_q_reg:Q oDFF_24_q_reg:D 32.9333
C1111 oDFF_29_q_reg:D 0 2.15531e-16
C1112 DFF_29_q_reg:Q 0 9.48687e-16
R984 DFF_29_q_reg:Q oDFF_29_q_reg:D 27.7333
C1113 oDFF_30_q_reg:D 0 2.58633e-16
C1114 DFF_30_q_reg:Q 0 7.29271e-16
R985 DFF_30_q_reg:Q oDFF_30_q_reg:D 27.7333
C1115 c0_U86:A 0 7.60586e-16
C1116 c0_U55:B 0 6.96951e-16
C1117 c0_U28:B 0 3.28473e-16
C1118 c0_U19:B 0 5.60475e-17
C1119 c0_U5:Y 0 1.20156e-15
C1120 c0_n5:7 0 1.31996e-15
R986 c0_U5:Y c0_n5:7 29.51
R987 c0_U5:Y c0_U86:A 37.3713
R988 c0_U5:Y c0_U55:B 29
R989 c0_U19:B c0_n5:7 6.4
R990 c0_U28:B c0_n5:7 23.6
R991 c0_U86:A c0_n5:7 82.1496
C1121 c0_U144:B 0 7.90441e-16
C1122 c0_U20:A 0 6.52534e-16
C1123 c0_U15:Y 0 4.15484e-16
R992 c0_U15:Y c0_U20:A 43.3783
R993 c0_U15:Y c0_U144:B 45.8689
R994 c0_U20:A c0_U144:B 42.2317
C1124 c0_U21:Y 0 8.99393e-16
C1125 c0_U20:B 0 6.89254e-16
R995 c0_U21:Y c0_U20:B 32.3333
C1126 c0_U32:Y 0 6.48392e-16
C1127 c0_U31:B 0 8.65042e-16
R996 c0_U32:Y c0_U31:B 32.2
C1128 c0_U42:Y 0 8.62953e-16
C1129 c0_U41:B 0 4.42179e-16
R997 c0_U42:Y c0_U41:B 28.9333
C1130 c0_U49:Y 0 5.88914e-16
C1131 c0_U48:B 0 3.54358e-16
C1132 c0_n43:3 0 2.31953e-15
R998 c0_U49:Y c0_n43:3 9.93333
R999 c0_U48:B c0_n43:3 26.5333
C1133 c0_U56:Y 0 3.38039e-16
C1134 c0_U55:C 0 1.43055e-15
R1000 c0_U56:Y c0_U55:C 18
C1135 c0_U101:Y 0 4.102e-16
C1136 c0_U97:A 0 3.11654e-16
R1001 c0_U101:Y c0_U97:A 2.2
C1137 c0_U99:Y 0 5.99501e-16
C1138 c0_U98:B 0 1.13902e-15
C1139 c0_n81:3 0 1.56839e-15
R1002 c0_U99:Y c0_n81:3 42.4
R1003 c0_U98:B c0_n81:3 9.73333
C1140 c0_U107:Y 0 5.22631e-16
C1141 c0_U105:A 0 5.62296e-16
C1142 c0_n88:3 0 1.15466e-15
R1004 c0_U107:Y c0_n88:3 8.4
R1005 c0_U105:A c0_n88:3 41.6667
C1143 c0_U140:Y 0 1.2493e-16
C1144 c0_U138:A 0 7.62552e-16
C1145 c0_n119:2 0 3.45371e-15
R1006 c0_U140:Y c0_n119:2 26.6667
R1007 c0_U138:A c0_n119:2 8.06667
C1146 c0_U143:Y 0 6.32878e-16
C1147 c0_U142:B 0 1.90315e-15
C1148 c0_n123:3 0 1.01555e-15
R1008 c0_U143:Y c0_n123:3 37.8667
R1009 c0_U142:B c0_n123:3 12.7333
C1149 c0_U151:Y 0 8.89322e-16
C1150 c0_U147:A 0 3.7935e-16
C1151 c0_n124:3 0 2.24099e-15
R1010 c0_U151:Y c0_n124:3 8.93333
R1011 c0_U147:A c0_n124:3 27
C1152 c0_U164:Y 0 1.10421e-15
C1153 c0_U160:A 0 1.46935e-16
C1154 c0_n134:2 0 1.07983e-15
R1012 c0_U164:Y c0_n134:2 25.6
R1013 c0_U160:A c0_n134:2 9.06667
C1155 c0_U163:Y 0 3.8523e-16
C1156 c0_U161:A 0 1.8506e-16
C1157 c0_n136:2 0 1.87606e-15
C1158 c0_n136:3 0 1.85511e-15
R1014 c0_U163:Y c0_n136:2 16.3333
R1015 c0_U161:A c0_n136:3 12.4
R1016 c0_n136:2 c0_n136:3 27.5333
C1159 c0_U180:Y 0 1.37277e-16
C1160 c0_U178:A 0 1.60524e-16
C1161 c0_n149:2 0 3.02781e-15
R1017 c0_U180:Y c0_n149:2 29.8667
R1018 c0_U178:A c0_n149:2 7.06667
C1162 c0_U183:Y 0 3.30697e-16
C1163 c0_U182:B 0 6.86325e-16
R1019 c0_U183:Y c0_U182:B 27.8
C1164 c0_n70:10 c0_n67:14 1.64033e-16
C1165 c0_n70:10 c0_U116:B 3.72187e-17
C1166 c0_n70:10 c0_U10:A 8.60455e-16
C1167 c0_U9:A c0_U10:A 3.84224e-17
C1168 c0_U125:Y c0_n67:14 3.37236e-17
C1169 c0_U125:Y c0_U117:B 3.65317e-17
C1170 c0_U128:B c0_n70:10 3.69819e-17
C1171 c0_U128:B c0_n70:8 5.83584e-18
C1172 iDFF_15_q_reg:Q c0_n70:10 1.94741e-16
C1173 iDFF_15_q_reg:Q c0_n70:8 3.80649e-17
C1174 iDFF_15_q_reg:Q c0_U90:A 7.05404e-17
C1175 c0_n9:11 c0_n70:10 1.68356e-17
C1176 c0_n9:11 c0_n67:14 1.38191e-16
C1177 c0_n9:11 c0_U116:B 7.51965e-17
C1178 c0_U9:Y c0_n70:10 2.36816e-17
C1179 c0_U9:Y c0_U10:A 5.96041e-18
C1180 c0_U116:A c0_n70:10 3.24675e-17
C1181 c0_U116:A c0_n67:14 3.94353e-17
C1182 c0_U116:A c0_U116:B 2.68591e-17
C1183 c0_U116:A c0_U10:A 3.69294e-18
C1184 c0_U113:A c0_n70:10 4.5522e-17
C1185 c0_U113:A c0_U117:A 3.26647e-17
C1186 c0_U113:A c0_n67:14 1.57162e-18
C1187 c0_U113:A c0_U116:B 1.037e-16
C1188 c0_U113:A c0_U10:A 6.54089e-20
C1189 c0_n10:9 c0_n9:11 3.51456e-17
C1190 c0_n10:9 c0_U61:B 1.02312e-16
C1191 c0_n10:9 IN_N57:7 4.60854e-16
C1192 c0_n10:9 c0_U170:B 3.51991e-17
C1193 c0_U59:B c0_U61:B 1.807e-17
C1194 c0_U10:Y IN_N57:7 3.15454e-17
C1195 c0_U113:B c0_U115:B 1.28141e-17
C1196 c0_U113:B c0_U117:A 2.88879e-16
C1197 clk__L2_N2:89 Qout_N729:5 5.38706e-17
C1198 clk__L2_N2:89 Qout_N729 6.54539e-17
C1199 clk__L2_N2:81 N13:4 7.2789e-17
C1200 clk__L2_N2:81 iDFF_4_q_reg:D 1.10467e-18
C1201 clk__L2_N2:75 c0_n67:12 5.09006e-17
C1202 clk__L2_N2:52 IN_N57:7 1.75535e-17
C1203 clk__L2_N2:52 c0_U60:A 8.75585e-17
C1204 iDFF_2_q_reg:CLK c0_n67:12 8.74338e-19
C1205 DFF_15_q_reg:CLK c0_U60:A 1.00273e-17
C1206 oDFF_4_q_reg:CLK N13:4 1.82171e-17
C1207 oDFF_4_q_reg:CLK N13 6.00033e-17
C1208 DFF_1_q_reg:CLK N13:4 1.35736e-18
C1209 iDFF_7_q_reg:CLK Qout_N729 1.30286e-16
C1210 oDFF_6_q_reg:CLK c0_n67:12 1.13423e-16
C1211 oDFF_6_q_reg:CLK oDFF_6_q_reg:Q 4.75654e-19
C1212 DFF_7_q_reg:CLK Qout_N729:5 1.26132e-18
C1213 DFF_7_q_reg:CLK Qout_N729:5 6.79808e-17
C1214 N136:4 N21:4 2.26922e-15
C1215 N136:4 N21 1.60949e-16
C1216 N136:3 N21:4 7.41138e-18
C1217 N136:3 N21:3 1.34604e-16
C1218 N136 N21:4 4.53895e-17
C1219 c0_n74:12 c0_n70:10 8.43431e-16
C1220 c0_n74:12 c0_U117:A 6.52293e-17
C1221 c0_n74:12 c0_U9:A 3.26353e-19
C1222 c0_n74:12 c0_n67:14 4.08175e-17
C1223 c0_n74:12 c0_U116:B 3.21173e-19
C1224 c0_n74:12 c0_U10:A 6.54265e-17
C1225 c0_n74:10 c0_n67:12 4.40242e-17
C1226 c0_n74:5 c0_n67:10 3.32003e-17
C1227 c0_n74:5 c0_U118:Y 5.57949e-19
C1228 c0_n74:5 c0_U88:A 4.30443e-17
C1229 c0_U88:B c0_U88:A 2.34932e-16
C1230 c0_U90:B c0_n70:10 1.3196e-16
C1231 c0_U90:B c0_U9:A 2.00988e-18
C1232 c0_U90:B c0_U90:A 3.4977e-17
C1233 c0_U90:B c0_U10:A 5.9927e-16
C1234 c0_n68:11 c0_n98:3 1.05527e-15
C1235 c0_n68:11 N136:4 2.78338e-16
C1236 c0_n68:11 N136:3 3.10411e-17
C1237 c0_n68:11 iDFF_40_q_reg:D 1.2454e-19
C1238 c0_n68:10 c0_n98:3 7.48205e-16
C1239 c0_n68:10 c0_n74:7 6.1509e-17
C1240 c0_n68:10 c0_n74:5 1.25091e-15
C1241 c0_n68:10 c0_n67:10 9.63653e-16
C1242 c0_n68:10 c0_U78:A 8.74338e-19
C1243 c0_n68:10 c0_U118:Y 3.57434e-17
C1244 c0_n68:10 c0_U88:A 7.56192e-17
C1245 c0_U78:B c0_n67:10 9.88789e-18
C1246 c0_n30:15 IN_N21:6 7.2654e-16
C1247 c0_n30:15 c0_U81:A 1.47212e-16
C1248 c0_n30:15 c0_U135:B 7.8744e-19
C1249 c0_n30:15 iDFF_6_q_reg:Q 2.94552e-17
C1250 c0_n30:15 N21:3 1.24148e-16
C1251 c0_n30:15 iDFF_6_q_reg:D 2.77635e-17
C1252 c0_U94:A IN_N21:8 3.17345e-16
C1253 c0_U94:A iDFF_6_q_reg:Q 3.79733e-17
C1254 c0_U173:Y N21:3 1.78005e-16
C1255 c0_n62:16 c0_n30:10 7.19801e-16
C1256 c0_n62:16 c0_U7:A 8.67401e-19
C1257 c0_n62:15 c0_n68:6 1.67982e-16
C1258 c0_n62:11 c0_n30:15 2.884e-17
C1259 c0_n62:8 c0_n30:10 5.82146e-17
C1260 c0_n140:5 c0_U115:A 4.34334e-17
C1261 c0_n140:2 c0_n10:9 1.53714e-15
C1262 c0_n140:2 c0_U115:A 3.70283e-17
C1263 c0_n140:2 IN_N57:7 1.27104e-16
C1264 c0_n140:2 c0_U170:B 3.18486e-19
C1265 c0_n146:4 c0_n62:15 5.96581e-16
C1266 c0_n146:4 c0_n62:8 1.46447e-17
C1267 c0_n146:4 N21:4 4.75768e-16
C1268 c0_n146:4 N21:3 1.39234e-17
C1269 c0_U174:A N21:4 3.96722e-17
C1270 c0_U176:Y c0_n62:8 3.4235e-17
C1271 IN_N37:8 c0_n62:8 1.10511e-16
C1272 c0_U135:A c0_n62:8 1.42656e-16
C1273 c0_U135:A c0_U132:A 3.86076e-19
C1274 c0_n54:12 c0_n140:5 1.26646e-15
C1275 c0_n54:12 c0_U165:B 5.88054e-17
C1276 c0_n54:8 c0_n10:11 3.20991e-16
C1277 c0_n54:8 c0_U59:B 2.85287e-17
C1278 c0_n54:8 c0_U68:B 1.42426e-17
C1279 c0_n54:8 clk__L2_N2:52 2.75085e-16
C1280 c0_n54:8 iDFF_14_q_reg:CLK 1.84877e-17
C1281 c0_U66:Y c0_U165:B 9.00968e-17
C1282 c0_U59:A clk__L2_N2:52 1.95083e-18
C1283 c0_U61:A clk__L2_N2:52 1.35859e-16
C1284 c0_n59:6 c0_n54:12 3.38025e-18
C1285 c0_n59:6 c0_n54:8 4.01138e-16
C1286 c0_n59:6 c0_U65:A 9.91808e-17
C1287 c0_n59:6 c0_U63:A 1.25322e-16
C1288 c0_n59:6 c0_n10:11 4.10053e-17
C1289 c0_n59:6 c0_U68:B 1.1182e-16
C1290 c0_U70:A c0_n9:11 6.11075e-17
C1291 c0_U70:A c0_U70:B 1.80998e-16
C1292 c0_U70:A c0_U61:B 4.41226e-17
C1293 iDFF_10_q_reg:D c0_U72:A 1.51279e-16
C1294 iDFF_10_q_reg:D c0_U74:A 2.76662e-17
C1295 N134:6 N130:6 5.5486e-19
C1296 N134:6 N130:4 5.95178e-17
C1297 N134:3 N130:4 3.42693e-16
C1298 N134:3 N130 5.39357e-16
C1299 IN_N137:20 N134:6 3.86302e-17
C1300 IN_N137:20 N130:6 5.95573e-17
C1301 IN_N137:20 iDFF_34_q_reg:D 5.76238e-18
C1302 IN_N137:19 N134:6 4.08581e-17
C1303 IN_N137:19 N130:4 3.42261e-17
C1304 IN_N137:19 N129:4 5.28162e-17
C1305 IN_N137:19 iDFF_33_q_reg:D 2.92662e-18
C1306 IN_N137:16 N134:6 6.57947e-18
C1307 c0_U145:B c0_n68:6 3.21729e-16
C1308 c0_U110:B N130:6 2.50977e-16
C1309 c0_U124:B N134:6 4.13388e-17
C1310 c0_U124:B N130:4 4.72612e-17
C1311 c0_U124:B N129:4 2.8685e-16
C1312 iDFF_41_q_reg:Q N134:6 1.32148e-19
C1313 c0_n21:7 c0_n62:16 1.19163e-16
C1314 c0_n21:7 c0_n62:8 2.8589e-17
C1315 c0_n21:7 c0_U114:C 2.59086e-17
C1316 c0_n21:7 c0_n30:10 1.25968e-16
C1317 c0_n21:7 c0_U112:A 5.6834e-17
C1318 c0_n21:7 IN_N37:8 3.50951e-17
C1319 c0_n21:7 c0_U135:A 3.38106e-16
C1320 c0_U114:A c0_U8:A 5.75968e-17
C1321 c0_U114:A c0_U114:C 8.67401e-19
C1322 c0_U116:Y c0_n9:11 1.5953e-16
C1323 c0_n27:5 c0_U176:Y 5.975e-16
C1324 c0_n27:5 c0_n62:16 1.44345e-16
C1325 c0_n27:5 c0_n62:8 2.72531e-17
C1326 c0_n27:5 c0_U114:C 1.13521e-16
C1327 c0_n27:5 c0_n30:10 2.02005e-15
C1328 c0_n27:5 c0_U34:C 3.57434e-17
C1329 c0_n27:5 c0_n21:7 2.37765e-16
C1330 c0_U115:Y c0_U114:C 1.72879e-16
C1331 c0_U114:B c0_n62:16 3.86076e-19
C1332 c0_U114:B c0_U114:C 1.62084e-19
C1333 c0_U114:B c0_n21:7 1.64328e-18
C1334 c0_U52:A c0_n21:7 3.60211e-17
C1335 c0_n29:6 c0_n27:5 3.13727e-16
C1336 c0_n29:6 c0_U33:A 5.55354e-17
C1337 c0_n29:4 c0_U33:A 9.18775e-17
C1338 c0_n29:4 c0_U52:A 4.06747e-16
C1339 c0_n51:9 c0_n30:10 2.72709e-17
C1340 c0_n51:8 c0_n30:10 3.75187e-16
C1341 c0_n51:8 c0_U34:C 3.76302e-17
C1342 c0_n51:8 c0_n29:6 4.15541e-16
C1343 c0_n51:8 c0_n29:4 3.55504e-17
C1344 c0_n51:8 c0_U34:B 2.77806e-18
C1345 c0_U66:B c0_n30:10 1.22845e-19
C1346 c0_n52:8 c0_U66:Y 3.7977e-17
C1347 c0_n52:8 c0_U56:A 4.84802e-17
C1348 c0_U56:B c0_U56:A 1.26717e-16
C1349 c0_U95:C c0_U66:Y 8.71171e-17
C1350 c0_U95:C c0_n51:9 1.21127e-16
C1351 c0_U95:C c0_n51:8 7.05963e-18
C1352 c0_n65:5 c0_n51:9 6.63479e-17
C1353 c0_n65:5 c0_U85:C 4.75129e-16
C1354 c0_U111:Y c0_n62:15 3.89176e-17
C1355 c0_U111:Y c0_n62:8 6.96578e-17
C1356 c0_U85:B c0_U85:C 2.54468e-17
C1357 c0_n83:7 c0_n21:7 2.55418e-16
C1358 c0_n83:7 c0_U43:A 2.29109e-18
C1359 c0_n91:5 c0_n62:16 6.88282e-17
C1360 c0_n91:5 c0_n62:8 2.14764e-17
C1361 c0_n91:5 c0_U114:C 2.7571e-17
C1362 c0_n91:5 c0_n51:8 7.94219e-17
C1363 c0_n91:5 c0_n30:10 1.13913e-16
C1364 c0_n91:5 c0_U34:C 1.56186e-18
C1365 c0_n91:5 c0_n29:6 1.55926e-17
C1366 c0_n91:5 c0_n29:4 1.56186e-18
C1367 c0_U108:B c0_n65:5 3.16768e-16
C1368 c0_U108:B c0_n51:8 7.21928e-17
C1369 c0_U108:B c0_n29:6 9.09096e-19
C1370 c0_U108:B c0_n29:4 2.85557e-16
C1371 c0_U108:B c0_U52:B 3.86076e-19
C1372 c0_U168:B c0_n65:5 3.69819e-17
C1373 c0_n8:6 c0_n59:6 5.34316e-16
C1374 c0_n8:6 c0_U72:A 3.43967e-17
C1375 c0_n8:6 c0_U74:A 2.88089e-17
C1376 c0_n8:6 c0_n54:12 3.22761e-17
C1377 c0_n8:6 c0_U65:A 9.58657e-18
C1378 c0_n8:5 c0_n52:8 1.14472e-16
C1379 c0_n8:5 c0_U75:A 5.97566e-17
C1380 c0_U63:B c0_n59:6 1.02472e-17
C1381 c0_U63:B c0_U65:A 1.17895e-16
C1382 c0_U8:Y c0_n54:12 5.70568e-17
C1383 c0_U34:A c0_n52:8 7.05481e-17
C1384 c0_U72:B c0_U72:A 9.62061e-18
C1385 clk__L2_N1:85 c0_U72:A 4.55238e-17
C1386 clk__L2_N1:85 c0_U74:A 1.40325e-17
C1387 clk__L2_N1:85 c0_n8:6 7.88887e-17
C1388 clk__L2_N1:85 c0_U72:B 1.54182e-16
C1389 clk__L2_N1:85 N37:3 7.31226e-17
C1390 clk__L2_N1:85 iDFF_10_q_reg:D 4.62532e-17
C1391 clk__L2_N1:84 IN_N137:20 3.13332e-18
C1392 clk__L2_N1:84 c0_U145:B 8.8681e-17
C1393 clk__L2_N1:84 c0_U110:B 9.46502e-17
C1394 clk__L2_N1:84 N130:6 1.43313e-17
C1395 clk__L2_N1:84 iDFF_34_q_reg:D 5.61797e-19
C1396 clk__L2_N1:79 N37:3 7.44857e-18
C1397 clk__L2_N1:76 c0_U72:A 8.22866e-17
C1398 clk__L2_N1:76 c0_U75:Y 3.91908e-19
C1399 clk__L2_N1:76 c0_U75:A 1.26955e-16
C1400 clk__L2_N1:76 c0_n8:6 4.57852e-17
C1401 clk__L2_N1:76 c0_n8:5 4.24249e-17
C1402 clk__L2_N1:76 c0_U72:B 4.78207e-19
C1403 clk__L2_N1:76 iDFF_10_q_reg:D 2.62762e-17
C1404 clk__L2_N1:70 IN_N137:19 3.38783e-16
C1405 clk__L2_N1:70 IN_N137:16 8.89307e-17
C1406 clk__L2_N1:70 N134:6 4.14112e-17
C1407 clk__L2_N1:70 N130:6 1.48155e-17
C1408 clk__L2_N1:70 N130:4 3.37243e-17
C1409 clk__L2_N1:70 N129:4 8.99001e-19
C1410 clk__L2_N1:70 iDFF_33_q_reg:D 4.88516e-18
C1411 clk__L2_N1:64 N129:4 1.11898e-16
C1412 clk__L2_N1:64 N129 9.91248e-17
C1413 clk__L2_N1:64 N17:4 1.03751e-16
C1414 clk__L2_N1:64 iDFF_5_q_reg:D 1.09612e-17
C1415 clk__L2_I1:Y iDFF_38_q_reg:D 8.66868e-20
C1416 DFF_9_q_reg:CLK N37:3 5.13476e-17
C1417 DFF_10_q_reg:CLK iDFF_10_q_reg:D 2.68636e-19
C1418 oDFF_9_q_reg:CLK N37:3 2.76217e-17
C1419 oDFF_9_q_reg:CLK N37:2 5.82964e-17
C1420 iDFF_34_q_reg:CLK IN_N137:20 6.19574e-17
C1421 iDFF_34_q_reg:CLK c0_U110:B 8.52131e-19
C1422 iDFF_34_q_reg:CLK iDFF_34_q_reg:D 2.70915e-17
C1423 iDFF_34_q_reg:CLK IN_N137:20 1.88058e-18
C1424 iDFF_34_q_reg:CLK iDFF_34_q_reg:D 1.09519e-17
C1425 iDFF_38_q_reg:CLK c0_n52:8 4.82772e-17
C1426 iDFF_38_q_reg:CLK c0_U75:A 4.44133e-19
C1427 iDFF_38_q_reg:CLK c0_n27:5 3.79686e-17
C1428 iDFF_38_q_reg:CLK c0_U33:A 4.25315e-17
C1429 iDFF_38_q_reg:CLK c0_U52:A 6.97818e-17
C1430 iDFF_38_q_reg:CLK c0_n8:5 6.72928e-17
C1431 iDFF_38_q_reg:CLK c0_U34:A 9.48258e-18
C1432 iDFF_38_q_reg:CLK iDFF_38_q_reg:D 1.56924e-17
C1433 iDFF_13_q_reg:CLK c0_U8:Y 3.18914e-17
C1434 iDFF_40_q_reg:CLK N130:6 5.35766e-20
C1435 iDFF_33_q_reg:CLK IN_N137:19 5.07851e-19
C1436 iDFF_33_q_reg:CLK N130:4 3.86076e-19
C1437 iDFF_20_q_reg:CLK IN_N137:19 3.21173e-19
C1438 iDFF_20_q_reg:CLK IN_N137:16 3.86076e-19
C1439 iDFF_37_q_reg:CLK IN_N137:16 5.56164e-18
C1440 iDFF_36_q_reg:CLK c0_U124:B 2.12005e-18
C1441 iDFF_35_q_reg:CLK N17:4 1.24652e-17
C1442 iDFF_5_q_reg:CLK N17:4 1.3675e-18
C1443 iDFF_5_q_reg:CLK iDFF_5_q_reg:D 4.57307e-17
C1444 iDFF_41_q_reg:CLK N134:6 4.37169e-17
C1445 iDFF_41_q_reg:CLK N130:4 1.30374e-17
C1446 iDFF_41_q_reg:CLK N129:4 1.27084e-16
C1447 iDFF_41_q_reg:CLK N129 2.72491e-17
C1448 oDFF_5_q_reg:CLK N17:4 2.51102e-17
C1449 DFF_24_q_reg:CLK IN_N137:19 7.80704e-19
C1450 DFF_24_q_reg:CLK IN_N137:16 1.07905e-17
C1451 DFF_24_q_reg:CLK c0_U124:B 7.10178e-19
C1452 DFF_24_q_reg:CLK iDFF_41_q_reg:Q 3.84146e-18
C1453 clk__L1_N0:7 clk__L2_I1:Y 1.47119e-18
C1454 clk__L1_N0:7 clk__L2_I1:Y 1.3511e-17
C1455 clk__L1_N0:7 iDFF_34_q_reg:CLK 4.50133e-19
C1456 clk__L1_N0:7 iDFF_38_q_reg:CLK 3.90761e-17
C1457 clk__L1_N0:7 iDFF_38_q_reg:D 1.22394e-16
C1458 clk__L1_N0:6 IN_N137:20 3.64294e-17
C1459 clk__L1_N0:6 IN_N137:19 3.78325e-17
C1460 clk__L1_N0:6 IN_N137:16 1.51132e-16
C1461 clk__L1_N0:6 c0_U172:A 3.94319e-18
C1462 clk__L1_N0:6 c0_U159:B 3.29374e-17
C1463 clk__L1_N0:6 c0_U124:B 3.59969e-17
C1464 clk__L1_N0:6 iDFF_41_q_reg:Q 2.82744e-18
C1465 clk__L1_N0:6 clk__L2_N1:70 2.41855e-16
C1466 clk__L1_N0:6 iDFF_37_q_reg:CLK 1.36657e-17
C1467 clk__L1_N0:6 iDFF_41_q_reg:CLK 3.85308e-17
C1468 clk__L1_N0:6 DFF_24_q_reg:CLK 3.86702e-16
C1469 clk__L1_N0:6 N134:6 1.88002e-15
C1470 clk__L1_N0:6 iDFF_38_q_reg:D 6.05909e-17
C1471 clk__L1_I0:Y N134:6 2.86368e-19
C1472 clk__L2_I2:A c0_n70:8 1.07355e-16
C1473 clk__L2_I2:A c0_U80:A 9.88006e-19
C1474 clk__L2_I2:A c0_n62:15 4.09781e-17
C1475 clk__L2_I2:A c0_n62:11 4.5177e-17
C1476 clk__L2_I2:A c0_U133:Y 3.80067e-17
C1477 clk__L2_I2:A clk__L2_N2:75 6.09093e-16
C1478 clk__L2_I2:A iDFF_2_q_reg:CLK 1.2417e-18
C1479 clk__L2_I2:A clk__L2_I2:Y 5.57949e-19
C1480 clk__L2_I1:A clk__L2_I1:Y 2.98416e-18
C1481 c0_n41:11 c0_U108:B 1.53706e-17
C1482 c0_n41:11 iDFF_38_q_reg:CLK 3.03349e-16
C1483 c0_U52:Y c0_U108:B 2.17225e-16
C1484 c0_U52:Y iDFF_38_q_reg:CLK 1.50741e-17
C1485 c0_n103:6 c0_n146:4 1.04372e-16
C1486 c0_n103:6 c0_n68:6 7.77276e-18
C1487 c0_n103:6 c0_U85:Y 4.83428e-17
C1488 c0_n103:6 c0_n65:5 3.21173e-19
C1489 c0_n103:6 c0_U111:Y 1.01577e-16
C1490 c0_n103:5 c0_n146:4 1.59807e-16
C1491 c0_n103:5 c0_n68:6 4.8584e-17
C1492 c0_U122:B c0_n146:4 2.64297e-17
C1493 c0_n46:6 c0_n103:6 9.00393e-16
C1494 c0_n46:6 c0_U108:B 2.74326e-16
C1495 c0_n46:6 c0_U168:B 6.25685e-17
C1496 c0_n46:6 c0_n65:5 5.54285e-16
C1497 c0_U1:A c0_n65:5 1.22064e-17
C1498 c0_U53:A c0_n103:6 1.79046e-17
C1499 c0_n111:4 c0_n83:7 1.67012e-16
C1500 c0_n111:4 c0_n83:5 3.46456e-17
C1501 c0_n111:4 c0_n65:5 2.74502e-16
C1502 c0_n111:4 c0_U76:B 3.07386e-19
C1503 c0_n111:4 c0_U95:B 1.32442e-17
C1504 c0_n111:4 c0_n51:9 2.95547e-16
C1505 c0_n111:4 c0_U85:C 6.0595e-17
C1506 c0_n111:4 c0_n29:9 1.24731e-15
C1507 c0_n111:4 c0_n29:4 5.47321e-16
C1508 c0_n111:4 c0_U53:Y 3.69819e-17
C1509 c0_n111:4 c0_U52:B 1.29209e-19
C1510 c0_n111:4 c0_n21:7 5.14789e-16
C1511 c0_n111:4 c0_U43:A 5.84764e-17
C1512 c0_n111:4 clk__L2_I2:A 1.15505e-17
C1513 c0_n111:3 clk__L2_I2:A 3.61838e-16
C1514 c0_U137:B clk__L1_N0:7 1.07592e-18
C1515 c0_U137:B clk__L2_I2:A 2.69756e-17
C1516 c0_U137:B clk__L2_I1:A 5.46702e-17
C1517 c0_U129:B clk__L2_I2:A 2.69756e-17
C1518 N135:4 iDFF_23_q_reg:CLK 1.479e-16
C1519 N135:4 oDFF_24_q_reg:CLK 4.12764e-16
C1520 N135:4 iDFF_24_q_reg:CLK 3.57316e-17
C1521 c0_n32:14 c0_n103:6 1.56221e-16
C1522 c0_n32:14 c0_U53:A 1.24163e-16
C1523 c0_n32:9 c0_n51:8 5.32382e-18
C1524 c0_n32:9 c0_U56:A 6.34109e-17
C1525 c0_n32:9 c0_U86:Y 3.80838e-16
C1526 c0_U86:B c0_U86:Y 2.0451e-17
C1527 c0_U11:A c0_n51:8 2.6361e-17
C1528 c0_U36:A c0_n41:7 1.22212e-16
C1529 c0_U36:A c0_U45:B 3.4643e-17
C1530 c0_U104:Y c0_n103:6 1.63737e-16
C1531 iDFF_31_q_reg:D DFF_31_q_reg:CLK 7.47406e-19
C1532 iDFF_31_q_reg:D iDFF_31_q_reg:CLK 2.07412e-16
C1533 IN_N77:4 c0_n41:7 1.49852e-15
C1534 IN_N77:4 c0_U45:B 6.44755e-17
C1535 IN_N77:4 c0_U36:A 5.27092e-17
C1536 IN_N77:4 c0_U45:A 7.00395e-17
C1537 c0_U179:A c0_n41:7 3.22297e-17
C1538 IN_N81:12 clk__L1_N0:7 4.42503e-16
C1539 c0_U41:A clk__L1_N0:7 3.91481e-17
C1540 c0_U150:B clk__L1_N0:7 7.22252e-17
C1541 c0_n35:15 c0_n83:5 4.90634e-16
C1542 c0_n35:15 c0_U164:B 7.77227e-21
C1543 c0_n35:15 clk__L1_N0:7 7.33841e-17
C1544 c0_n35:14 c0_n83:5 6.53292e-17
C1545 c0_n35:14 clk__L1_N0:7 5.06557e-17
C1546 c0_n35:11 c0_U96:Y 2.70113e-16
C1547 c0_U5:A c0_n52:8 1.36803e-16
C1548 c0_U5:A c0_U96:Y 3.69819e-17
C1549 c0_U57:A clk__L1_N0:7 1.88481e-16
C1550 c0_U11:Y c0_n83:5 1.00012e-16
C1551 c0_U11:Y c0_U11:A 2.1968e-17
C1552 c0_U26:B c0_n32:9 8.69422e-17
C1553 c0_U26:B c0_U86:B 1.77973e-17
C1554 c0_U26:B IN_N125:6 5.61167e-18
C1555 c0_U26:B c0_U106:A 2.42359e-16
C1556 c0_U17:B IN_N125:6 1.66991e-18
C1557 c0_U96:A c0_U86:B 8.66868e-20
C1558 c0_U96:A IN_N125:6 4.50133e-19
C1559 c0_U11:Y c0_n32:9 2.35473e-16
C1560 c0_U11:Y c0_U11:A 4.09762e-16
C1561 c0_U11:Y c0_U106:A 3.56814e-16
C1562 c0_n17:13 c0_n52:8 6.53946e-17
C1563 c0_n17:13 c0_U96:Y 2.12005e-18
C1564 c0_n17:13 c0_U56:B 1.25377e-16
C1565 c0_n17:13 c0_U56:A 1.24629e-16
C1566 c0_n17:13 c0_U86:Y 2.22941e-17
C1567 c0_n17:13 c0_U26:B 1.52983e-16
C1568 c0_n17:13 c0_U17:B 1.31561e-17
C1569 c0_n17:13 c0_U96:A 4.11693e-16
C1570 c0_U24:Y c0_n52:8 3.45541e-16
C1571 c0_U24:Y c0_U56:B 3.09394e-17
C1572 c0_U24:Y c0_n51:8 8.46565e-16
C1573 c0_U24:Y c0_U56:A 5.28281e-17
C1574 c0_U24:Y c0_U11:Y 2.15429e-17
C1575 c0_n33:15 c0_n83:5 4.36539e-18
C1576 c0_n33:15 c0_n41:7 8.56773e-16
C1577 c0_n33:15 c0_U47:B 5.34252e-17
C1578 c0_n33:15 c0_U38:A 2.12097e-17
C1579 c0_n33:15 c0_U97:Y 1.30541e-18
C1580 c0_n33:15 c0_U47:A 5.72208e-17
C1581 c0_n33:15 c0_U97:Y 1.31895e-18
C1582 c0_n33:10 c0_n83:5 1.90907e-16
C1583 c0_n33:10 c0_U164:B 1.47228e-19
C1584 c0_n33:10 c0_n35:14 5.97261e-17
C1585 c0_n33:10 c0_U97:Y 2.10334e-18
C1586 c0_n33:10 c0_U11:Y 1.75576e-17
C1587 c0_U36:B c0_n41:7 4.83011e-16
C1588 c0_U36:B N135:4 1.26802e-16
C1589 c0_U43:Y c0_n83:5 6.16412e-17
C1590 c0_U43:Y c0_n35:15 4.12717e-17
C1591 c0_U43:Y c0_U11:Y 1.04641e-16
C1592 c0_U42:B c0_n83:5 1.47228e-19
C1593 c0_U40:B c0_U47:B 9.21312e-17
C1594 c0_U38:B c0_U47:A 1.58257e-17
C1595 c0_n37:16 c0_U51:B 2.73363e-19
C1596 c0_n37:16 c0_U49:B 1.19089e-17
C1597 c0_n37:13 c0_n111:4 5.32485e-16
C1598 c0_n37:13 c0_n35:15 6.14968e-16
C1599 c0_n37:13 c0_U11:Y 2.79996e-16
C1600 c0_n37:13 c0_U55:A 3.76302e-17
C1601 c0_U56:C c0_n35:15 2.88796e-17
C1602 c0_U12:A c0_U138:Y 6.10821e-17
C1603 c0_U12:A c0_U55:A 6.63887e-17
C1604 c0_U49:A c0_U49:B 1.75619e-16
C1605 c0_n39:14 c0_n65:6 3.57826e-16
C1606 c0_n39:14 c0_U76:B 2.54468e-17
C1607 c0_n39:14 c0_n46:7 1.29139e-16
C1608 c0_n39:14 c0_U43:Y 4.37968e-16
C1609 c0_n39:14 c0_n29:9 2.75043e-17
C1610 c0_n39:14 c0_U53:Y 3.09478e-17
C1611 c0_n39:11 c0_n83:5 3.73236e-16
C1612 c0_n39:11 c0_U164:B 1.64328e-18
C1613 c0_n39:11 c0_n35:15 9.01866e-17
C1614 c0_n39:11 c0_n35:14 2.93034e-16
C1615 c0_n39:11 c0_U97:Y 3.68075e-17
C1616 c0_n39:11 c0_n33:10 1.60999e-16
C1617 c0_n39:11 c0_U42:B 3.86076e-19
C1618 c0_n39:11 clk__L1_N0:7 4.48743e-16
C1619 c0_U54:A c0_n83:5 5.23332e-17
C1620 c0_U54:A c0_n46:7 2.28289e-16
C1621 c0_U54:A c0_n35:15 1.51052e-16
C1622 c0_U54:A c0_n33:10 1.89917e-18
C1623 c0_U54:A c0_U43:Y 1.72106e-17
C1624 c0_U54:A c0_U53:Y 9.05322e-17
C1625 c0_U76:C c0_n29:9 1.39487e-19
C1626 c0_U51:A clk__L1_N0:7 3.29653e-17
C1627 c0_U42:A c0_n35:14 4.63945e-20
C1628 c0_U42:A c0_n33:10 2.68636e-19
C1629 c0_U42:A clk__L1_N0:7 1.62084e-19
C1630 c0_U147:Y clk__L1_N0:7 1.62022e-17
C1631 IN_N109:6 c0_n52:8 6.08767e-16
C1632 IN_N109:6 c0_U96:Y 3.42759e-17
C1633 c0_U106:B c0_n52:8 2.12888e-17
C1634 c0_n23:9 c0_n52:8 5.6575e-17
C1635 c0_n23:9 c0_U96:Y 2.5314e-17
C1636 c0_n23:9 c0_U56:A 2.35114e-17
C1637 c0_n23:9 c0_U86:Y 3.33051e-19
C1638 c0_n23:9 c0_n17:13 2.97126e-17
C1639 c0_n23:9 c0_n17:9 3.21173e-19
C1640 c0_n23:9 c0_U24:Y 3.55504e-17
C1641 c0_n23:9 c0_U26:B 1.86686e-16
C1642 c0_n23:9 c0_U96:A 5.67696e-19
C1643 c0_n23:9 c0_U11:Y 2.34097e-17
C1644 c0_n23:9 IN_N109:6 2.09769e-15
C1645 c0_n23:9 c0_U106:B 1.90092e-16
C1646 c0_n23:9 c0_U139:B 3.19157e-17
C1647 c0_n23:7 c0_n52:8 5.21814e-16
C1648 c0_n23:7 c0_n51:8 1.64207e-16
C1649 c0_n23:7 c0_U24:Y 2.01188e-16
C1650 c0_n23:7 c0_U106:B 2.37978e-17
C1651 c0_U26:A IN_N109:6 2.83488e-17
C1652 c0_U28:A c0_n17:9 7.33009e-19
C1653 c0_U33:Y c0_n52:8 4.73301e-18
C1654 c0_U33:Y c0_n51:8 2.06459e-17
C1655 c0_U32:A c0_n17:9 2.55205e-17
C1656 c0_U32:A c0_U21:A 8.9745e-19
C1657 c0_n12:8 c0_n111:4 1.49041e-15
C1658 c0_n12:8 c0_U138:Y 6.63122e-17
C1659 c0_n12:8 c0_n83:7 9.19899e-17
C1660 c0_n12:8 c0_n83:5 4.29235e-17
C1661 c0_n12:8 c0_n39:14 1.52542e-18
C1662 c0_n12:8 c0_U76:C 6.093e-17
C1663 c0_n12:7 c0_U28:A 3.11988e-16
C1664 c0_n12:7 c0_U32:A 1.9623e-16
C1665 c0_n12:7 c0_n17:9 2.84915e-17
C1666 c0_n12:7 c0_U21:A 6.19269e-16
C1667 c0_U21:B c0_U21:A 1.95104e-16
C1668 c0_U76:A c0_n111:4 3.43035e-17
C1669 c0_U76:A c0_n39:14 6.22983e-17
C1670 c0_U30:B c0_U28:A 1.32442e-17
C1671 c0_U149:A iDFF_21_q_reg:Q 5.74243e-17
C1672 c0_U14:A IN_N81:8 1.47228e-19
C1673 c0_U14:A iDFF_21_q_reg:Q 1.56749e-16
C1674 c0_U14:A iDFF_21_q_reg:Q 1.33293e-17
C1675 IN_N97:5 c0_U12:A 5.98433e-17
C1676 IN_N97:5 c0_U160:Y 1.20329e-18
C1677 c0_U150:A c0_n37:16 7.53129e-17
C1678 c0_U150:A c0_U160:Y 1.88852e-17
C1679 c0_U150:A IN_N81:12 4.22035e-17
C1680 c0_U150:A c0_U41:A 9.13671e-17
C1681 clk__L2_N0:84 IN_N65:6 1.48872e-16
C1682 clk__L2_N0:84 iDFF_17_q_reg:Q 1.99643e-17
C1683 clk__L2_N0:84 N81:4 3.38871e-16
C1684 clk__L2_N0:73 IN_N97:7 1.01281e-16
C1685 clk__L2_N0:66 iDFF_27_q_reg:D 7.44857e-18
C1686 iDFF_21_q_reg:CLK N81:4 8.4988e-18
C1687 DFF_17_q_reg:CLK N81:4 5.07851e-19
C1688 iDFF_39_q_reg:CLK c0_U38:A 1.89552e-16
C1689 iDFF_39_q_reg:CLK c0_U47:A 5.47918e-17
C1690 iDFF_39_q_reg:CLK c0_n33:15 1.10133e-16
C1691 iDFF_39_q_reg:CLK c0_U38:B 6.53696e-18
C1692 iDFF_39_q_reg:CLK c0_U14:A 3.96716e-17
C1693 clk__L2_I0:Y iDFF_25_q_reg:Q 1.93923e-17
C1694 DFF_30_q_reg:CLK IN_N97:7 1.90026e-17
C1695 iDFF_27_q_reg:CLK iDFF_27_q_reg:D 1.61632e-17
C1696 iDFF_28_q_reg:CLK iDFF_27_q_reg:D 1.03405e-16
C1697 DFF_21_q_reg:CLK clk__L1_N0:7 3.24569e-16
C1698 DFF_21_q_reg:CLK clk__L2_I0:A 3.76302e-17
C1699 oDFF_17_q_reg:CLK N81:4 3.21173e-19
Xclk__L2_I2 clk__L2_I2:A clk__L2_I2:gnd clk__L2_I2:Y clk__L2_I2:vdd INVX8
Xclk__L2_I1 clk__L2_I1:A clk__L2_I1:gnd clk__L2_I1:Y clk__L2_I1:vdd INVX8
Xclk__L2_I0 clk__L2_I0:A clk__L2_I0:gnd clk__L2_I0:Y clk__L2_I0:vdd INVX8
Xclk__L1_I0 clk__L1_I0:A clk__L1_I0:gnd clk__L1_I0:Y clk__L1_I0:vdd INVX8
Xc0_U1 c0_U1:A c0_U1:gnd c0_U1:Y c0_U1:vdd INVX2
Xc0_U2 c0_U2:A c0_U2:gnd c0_U2:Y c0_U2:vdd INVX2
Xc0_U3 c0_U3:A c0_U3:gnd c0_U3:Y c0_U3:vdd INVX2
Xc0_U4 c0_U4:A c0_U4:gnd c0_U4:Y c0_U4:vdd INVX2
Xc0_U5 c0_U5:A c0_U5:gnd c0_U5:Y c0_U5:vdd INVX2
Xc0_U6 c0_U6:A c0_U6:gnd c0_U6:Y c0_U6:vdd INVX2
Xc0_U7 c0_U7:A c0_U7:gnd c0_U7:Y c0_U7:vdd INVX2
Xc0_U8 c0_U8:A c0_U8:gnd c0_U8:Y c0_U8:vdd INVX2
Xc0_U9 c0_U9:A c0_U9:gnd c0_U9:Y c0_U9:vdd INVX2
Xc0_U10 c0_U10:A c0_U10:gnd c0_U10:Y c0_U10:vdd INVX2
Xc0_U11 c0_U11:A c0_U11:gnd c0_U11:Y c0_U11:vdd INVX2
Xc0_U12 c0_U12:A c0_U12:gnd c0_U12:Y c0_U12:vdd INVX2
Xc0_U13 c0_U13:A c0_U13:gnd c0_U13:Y c0_U13:vdd INVX2
Xc0_U14 c0_U14:A c0_U14:gnd c0_U14:Y c0_U14:vdd INVX2
Xc0_U15 c0_U15:A c0_U15:gnd c0_U15:Y c0_U15:vdd INVX2
Xc0_U16 c0_U16:A c0_U16:B c0_U16:gnd c0_U16:Y c0_U16:vdd XNOR2X1
Xc0_U17 c0_U17:A c0_U17:B c0_U17:gnd c0_U17:Y c0_U17:vdd NAND2X1
Xc0_U18 c0_U18:A c0_U18:B c0_U18:gnd c0_U18:Y c0_U18:vdd XNOR2X1
Xc0_U19 c0_U19:A c0_U19:B c0_U19:gnd c0_U19:Y c0_U19:vdd NAND2X1
Xc0_U20 c0_U20:A c0_U20:B c0_U20:gnd c0_U20:Y c0_U20:vdd XOR2X1
Xc0_U21 c0_U21:A c0_U21:B c0_U21:gnd c0_U21:Y c0_U21:vdd NAND2X1
Xc0_U22 c0_U22:A c0_U22:B c0_U22:gnd c0_U22:Y c0_U22:vdd XNOR2X1
Xc0_U23 c0_U23:A c0_U23:B c0_U23:gnd c0_U23:Y c0_U23:vdd NAND2X1
Xc0_U24 c0_U24:A c0_U24:B c0_U24:gnd c0_U24:Y c0_U24:vdd AND2X1
Xc0_U25 c0_U25:A c0_U25:B c0_U25:gnd c0_U25:Y c0_U25:vdd XNOR2X1
Xc0_U26 c0_U26:A c0_U26:B c0_U26:gnd c0_U26:Y c0_U26:vdd NAND2X1
Xc0_U27 c0_U27:A c0_U27:B c0_U27:gnd c0_U27:Y c0_U27:vdd XNOR2X1
Xc0_U28 c0_U28:A c0_U28:B c0_U28:gnd c0_U28:Y c0_U28:vdd NAND2X1
Xc0_U29 c0_U29:A c0_U29:B c0_U29:gnd c0_U29:Y c0_U29:vdd XNOR2X1
Xc0_U30 c0_U30:A c0_U30:B c0_U30:gnd c0_U30:Y c0_U30:vdd NAND2X1
Xc0_U31 c0_U31:A c0_U31:B c0_U31:gnd c0_U31:Y c0_U31:vdd XNOR2X1
Xc0_U32 c0_U32:A c0_U32:B c0_U32:gnd c0_U32:Y c0_U32:vdd NAND2X1
Xc0_U33 c0_U33:A c0_U33:B c0_U33:gnd c0_U33:Y c0_U33:vdd AND2X1
Xc0_U34 c0_U34:A c0_U34:B c0_U34:C c0_U34:gnd c0_U34:Y c0_U34:vdd NAND3X1
Xc0_U35 c0_U35:A c0_U35:B c0_U35:gnd c0_U35:Y c0_U35:vdd XOR2X1
Xc0_U36 c0_U36:A c0_U36:B c0_U36:gnd c0_U36:Y c0_U36:vdd NOR2X1
Xc0_U37 c0_U37:A c0_U37:B c0_U37:gnd c0_U37:Y c0_U37:vdd XOR2X1
Xc0_U38 c0_U38:A c0_U38:B c0_U38:gnd c0_U38:Y c0_U38:vdd NOR2X1
Xc0_U39 c0_U39:A c0_U39:B c0_U39:gnd c0_U39:Y c0_U39:vdd XOR2X1
Xc0_U40 c0_U40:A c0_U40:B c0_U40:gnd c0_U40:Y c0_U40:vdd NOR2X1
Xc0_U41 c0_U41:A c0_U41:B c0_U41:gnd c0_U41:Y c0_U41:vdd XOR2X1
Xc0_U42 c0_U42:A c0_U42:B c0_U42:gnd c0_U42:Y c0_U42:vdd NOR2X1
Xc0_U43 c0_U43:A c0_U43:B c0_U43:C c0_U43:gnd c0_U43:Y c0_U43:vdd NAND3X1
Xc0_U44 c0_U44:A c0_U44:B c0_U44:gnd c0_U44:Y c0_U44:vdd XOR2X1
Xc0_U45 c0_U45:A c0_U45:B c0_U45:gnd c0_U45:Y c0_U45:vdd NOR2X1
Xc0_U46 c0_U46:A c0_U46:B c0_U46:gnd c0_U46:Y c0_U46:vdd XOR2X1
Xc0_U47 c0_U47:A c0_U47:B c0_U47:gnd c0_U47:Y c0_U47:vdd NOR2X1
Xc0_U48 c0_U48:A c0_U48:B c0_U48:gnd c0_U48:Y c0_U48:vdd XOR2X1
Xc0_U49 c0_U49:A c0_U49:B c0_U49:gnd c0_U49:Y c0_U49:vdd NOR2X1
Xc0_U50 c0_U50:A c0_U50:B c0_U50:gnd c0_U50:Y c0_U50:vdd XOR2X1
Xc0_U51 c0_U51:A c0_U51:B c0_U51:gnd c0_U51:Y c0_U51:vdd NOR2X1
Xc0_U52 c0_U52:A c0_U52:B c0_U52:C c0_U52:gnd c0_U52:Y c0_U52:vdd NAND3X1
Xc0_U53 c0_U53:A c0_U53:B c0_U53:C c0_U53:gnd c0_U53:Y c0_U53:vdd OAI21X1
Xc0_U54 c0_U54:A c0_U54:B c0_U54:gnd c0_U54:Y c0_U54:vdd NAND2X1
Xc0_U55 c0_U55:A c0_U55:B c0_U55:C c0_U55:gnd c0_U55:Y c0_U55:vdd OAI21X1
Xc0_U56 c0_U56:A c0_U56:B c0_U56:C c0_U56:gnd c0_U56:Y c0_U56:vdd OAI21X1
Xc0_U57 c0_U57:A c0_U57:B c0_U57:gnd c0_U57:Y c0_U57:vdd NAND2X1
Xc0_U58 c0_U58:A c0_U58:B c0_U58:gnd c0_U58:Y c0_U58:vdd XNOR2X1
Xc0_U59 c0_U59:A c0_U59:B c0_U59:gnd c0_U59:Y c0_U59:vdd NAND2X1
Xc0_U60 c0_U60:A c0_U60:B c0_U60:gnd c0_U60:Y c0_U60:vdd XNOR2X1
Xc0_U61 c0_U61:A c0_U61:B c0_U61:gnd c0_U61:Y c0_U61:vdd NAND2X1
Xc0_U62 c0_U62:A c0_U62:B c0_U62:gnd c0_U62:Y c0_U62:vdd XNOR2X1
Xc0_U63 c0_U63:A c0_U63:B c0_U63:gnd c0_U63:Y c0_U63:vdd NAND2X1
Xc0_U64 c0_U64:A c0_U64:B c0_U64:gnd c0_U64:Y c0_U64:vdd XOR2X1
Xc0_U65 c0_U65:A c0_U65:B c0_U65:gnd c0_U65:Y c0_U65:vdd NAND2X1
Xc0_U66 c0_U66:A c0_U66:B c0_U66:gnd c0_U66:Y c0_U66:vdd AND2X1
Xc0_U67 c0_U67:A c0_U67:B c0_U67:gnd c0_U67:Y c0_U67:vdd XNOR2X1
Xc0_U68 c0_U68:A c0_U68:B c0_U68:gnd c0_U68:Y c0_U68:vdd NAND2X1
Xc0_U69 c0_U69:A c0_U69:B c0_U69:gnd c0_U69:Y c0_U69:vdd XNOR2X1
Xc0_U70 c0_U70:A c0_U70:B c0_U70:gnd c0_U70:Y c0_U70:vdd NAND2X1
Xc0_U71 c0_U71:A c0_U71:B c0_U71:gnd c0_U71:Y c0_U71:vdd XNOR2X1
Xc0_U72 c0_U72:A c0_U72:B c0_U72:gnd c0_U72:Y c0_U72:vdd NAND2X1
Xc0_U73 c0_U73:A c0_U73:B c0_U73:gnd c0_U73:Y c0_U73:vdd XNOR2X1
Xc0_U74 c0_U74:A c0_U74:B c0_U74:gnd c0_U74:Y c0_U74:vdd NAND2X1
Xc0_U75 c0_U75:A c0_U75:B c0_U75:gnd c0_U75:Y c0_U75:vdd AND2X1
Xc0_U76 c0_U76:A c0_U76:B c0_U76:C c0_U76:gnd c0_U76:Y c0_U76:vdd NAND3X1
Xc0_U77 c0_U77:A c0_U77:B c0_U77:gnd c0_U77:Y c0_U77:vdd XOR2X1
Xc0_U78 c0_U78:A c0_U78:B c0_U78:gnd c0_U78:Y c0_U78:vdd NOR2X1
Xc0_U79 c0_U79:A c0_U79:B c0_U79:gnd c0_U79:Y c0_U79:vdd XOR2X1
Xc0_U80 c0_U80:A c0_U80:B c0_U80:gnd c0_U80:Y c0_U80:vdd NOR2X1
Xc0_U81 c0_U81:A c0_U81:B c0_U81:gnd c0_U81:Y c0_U81:vdd XOR2X1
Xc0_U82 c0_U82:A c0_U82:B c0_U82:gnd c0_U82:Y c0_U82:vdd NOR2X1
Xc0_U83 c0_U83:A c0_U83:B c0_U83:gnd c0_U83:Y c0_U83:vdd XOR2X1
Xc0_U84 c0_U84:A c0_U84:B c0_U84:gnd c0_U84:Y c0_U84:vdd NOR2X1
Xc0_U85 c0_U85:A c0_U85:B c0_U85:C c0_U85:gnd c0_U85:Y c0_U85:vdd NAND3X1
Xc0_U86 c0_U86:A c0_U86:B c0_U86:gnd c0_U86:Y c0_U86:vdd NOR2X1
Xc0_U87 c0_U87:A c0_U87:B c0_U87:gnd c0_U87:Y c0_U87:vdd XOR2X1
Xc0_U88 c0_U88:A c0_U88:B c0_U88:gnd c0_U88:Y c0_U88:vdd NOR2X1
Xc0_U89 c0_U89:A c0_U89:B c0_U89:gnd c0_U89:Y c0_U89:vdd XOR2X1
Xc0_U90 c0_U90:A c0_U90:B c0_U90:gnd c0_U90:Y c0_U90:vdd NOR2X1
Xc0_U91 c0_U91:A c0_U91:B c0_U91:gnd c0_U91:Y c0_U91:vdd XOR2X1
Xc0_U92 c0_U92:A c0_U92:B c0_U92:gnd c0_U92:Y c0_U92:vdd NOR2X1
Xc0_U93 c0_U93:A c0_U93:B c0_U93:gnd c0_U93:Y c0_U93:vdd XOR2X1
Xc0_U94 c0_U94:A c0_U94:B c0_U94:gnd c0_U94:Y c0_U94:vdd NOR2X1
Xc0_U95 c0_U95:A c0_U95:B c0_U95:C c0_U95:gnd c0_U95:Y c0_U95:vdd NAND3X1
Xc0_U96 c0_U96:A c0_U96:B c0_U96:gnd c0_U96:Y c0_U96:vdd NOR2X1
Xc0_U97 c0_U97:A c0_U97:B c0_U97:gnd c0_U97:Y c0_U97:vdd XOR2X1
Xc0_U98 c0_U98:A c0_U98:B c0_U98:gnd c0_U98:Y c0_U98:vdd XOR2X1
Xc0_U99 c0_U99:A c0_U99:B c0_U99:gnd c0_U99:Y c0_U99:vdd XOR2X1
Xc0_U100 c0_U100:A c0_U100:B c0_U100:gnd c0_U100:Y c0_U100:vdd XOR2X1
Xc0_U101 c0_U101:A c0_U101:B c0_U101:gnd c0_U101:Y c0_U101:vdd XOR2X1
Xc0_U102 c0_U102:A c0_U102:B c0_U102:gnd c0_U102:Y c0_U102:vdd XOR2X1
Xc0_U103 c0_U103:A c0_U103:B c0_U103:gnd c0_U103:Y c0_U103:vdd NAND2X1
Xc0_U104 c0_U104:A c0_U104:B c0_U104:gnd c0_U104:Y c0_U104:vdd XOR2X1
Xc0_U105 c0_U105:A c0_U105:B c0_U105:gnd c0_U105:Y c0_U105:vdd XOR2X1
Xc0_U106 c0_U106:A c0_U106:B c0_U106:gnd c0_U106:Y c0_U106:vdd XOR2X1
Xc0_U107 c0_U107:A c0_U107:B c0_U107:gnd c0_U107:Y c0_U107:vdd XOR2X1
Xc0_U108 c0_U108:A c0_U108:B c0_U108:gnd c0_U108:Y c0_U108:vdd XOR2X1
Xc0_U109 c0_U109:A c0_U109:B c0_U109:gnd c0_U109:Y c0_U109:vdd XOR2X1
Xc0_U110 c0_U110:A c0_U110:B c0_U110:gnd c0_U110:Y c0_U110:vdd NAND2X1
Xc0_U111 c0_U111:A c0_U111:B c0_U111:C c0_U111:gnd c0_U111:Y c0_U111:vdd OAI21X1
Xc0_U112 c0_U112:A c0_U112:B c0_U112:gnd c0_U112:Y c0_U112:vdd NAND2X1
Xc0_U113 c0_U113:A c0_U113:B c0_U113:C c0_U113:gnd c0_U113:Y c0_U113:vdd OAI21X1
Xc0_U114 c0_U114:A c0_U114:B c0_U114:C c0_U114:gnd c0_U114:Y c0_U114:vdd OAI21X1
Xc0_U115 c0_U115:A c0_U115:B c0_U115:gnd c0_U115:Y c0_U115:vdd NOR2X1
Xc0_U116 c0_U116:A c0_U116:B c0_U116:gnd c0_U116:Y c0_U116:vdd NOR2X1
Xc0_U117 c0_U117:A c0_U117:B c0_U117:gnd c0_U117:Y c0_U117:vdd NAND2X1
Xc0_U118 c0_U118:A c0_U118:B c0_U118:gnd c0_U118:Y c0_U118:vdd XOR2X1
Xc0_U119 c0_U119:A c0_U119:B c0_U119:gnd c0_U119:Y c0_U119:vdd XOR2X1
Xc0_U120 c0_U120:A c0_U120:B c0_U120:gnd c0_U120:Y c0_U120:vdd XOR2X1
Xc0_U121 c0_U121:A c0_U121:B c0_U121:gnd c0_U121:Y c0_U121:vdd XOR2X1
Xc0_U122 c0_U122:A c0_U122:B c0_U122:gnd c0_U122:Y c0_U122:vdd XOR2X1
Xc0_U123 c0_U123:A c0_U123:B c0_U123:gnd c0_U123:Y c0_U123:vdd XOR2X1
Xc0_U124 c0_U124:A c0_U124:B c0_U124:gnd c0_U124:Y c0_U124:vdd NAND2X1
Xc0_U125 c0_U125:A c0_U125:B c0_U125:gnd c0_U125:Y c0_U125:vdd XOR2X1
Xc0_U126 c0_U126:A c0_U126:B c0_U126:gnd c0_U126:Y c0_U126:vdd XOR2X1
Xc0_U127 c0_U127:A c0_U127:B c0_U127:gnd c0_U127:Y c0_U127:vdd XOR2X1
Xc0_U128 c0_U128:A c0_U128:B c0_U128:gnd c0_U128:Y c0_U128:vdd XOR2X1
Xc0_U129 c0_U129:A c0_U129:B c0_U129:gnd c0_U129:Y c0_U129:vdd XOR2X1
Xc0_U130 c0_U130:A c0_U130:B c0_U130:gnd c0_U130:Y c0_U130:vdd XOR2X1
Xc0_U131 c0_U131:A c0_U131:B c0_U131:gnd c0_U131:Y c0_U131:vdd NAND2X1
Xc0_U132 c0_U132:A c0_U132:B c0_U132:gnd c0_U132:Y c0_U132:vdd NAND2X1
Xc0_U133 c0_U133:A c0_U133:B c0_U133:gnd c0_U133:Y c0_U133:vdd XOR2X1
Xc0_U134 c0_U134:A c0_U134:B c0_U134:gnd c0_U134:Y c0_U134:vdd XOR2X1
Xc0_U135 c0_U135:A c0_U135:B c0_U135:gnd c0_U135:Y c0_U135:vdd XOR2X1
Xc0_U136 c0_U136:A c0_U136:B c0_U136:gnd c0_U136:Y c0_U136:vdd XOR2X1
Xc0_U137 c0_U137:A c0_U137:B c0_U137:gnd c0_U137:Y c0_U137:vdd XOR2X1
Xc0_U138 c0_U138:A c0_U138:B c0_U138:gnd c0_U138:Y c0_U138:vdd XNOR2X1
Xc0_U139 c0_U139:A c0_U139:B c0_U139:gnd c0_U139:Y c0_U139:vdd XOR2X1
Xc0_U140 c0_U140:A c0_U140:B c0_U140:gnd c0_U140:Y c0_U140:vdd XNOR2X1
Xc0_U141 c0_U141:A c0_U141:B c0_U141:gnd c0_U141:Y c0_U141:vdd XOR2X1
Xc0_U142 c0_U142:A c0_U142:B c0_U142:gnd c0_U142:Y c0_U142:vdd XNOR2X1
Xc0_U143 c0_U143:A c0_U143:B c0_U143:gnd c0_U143:Y c0_U143:vdd XOR2X1
Xc0_U144 c0_U144:A c0_U144:B c0_U144:gnd c0_U144:Y c0_U144:vdd XOR2X1
Xc0_U145 c0_U145:A c0_U145:B c0_U145:gnd c0_U145:Y c0_U145:vdd NAND2X1
Xc0_U146 c0_U146:A c0_U146:B c0_U146:gnd c0_U146:Y c0_U146:vdd NAND2X1
Xc0_U147 c0_U147:A c0_U147:B c0_U147:gnd c0_U147:Y c0_U147:vdd XOR2X1
Xc0_U148 c0_U148:A c0_U148:B c0_U148:gnd c0_U148:Y c0_U148:vdd XOR2X1
Xc0_U149 c0_U149:A c0_U149:B c0_U149:gnd c0_U149:Y c0_U149:vdd XOR2X1
Xc0_U150 c0_U150:A c0_U150:B c0_U150:gnd c0_U150:Y c0_U150:vdd XOR2X1
Xc0_U151 c0_U151:A c0_U151:B c0_U151:gnd c0_U151:Y c0_U151:vdd XOR2X1
Xc0_U152 c0_U152:A c0_U152:B c0_U152:gnd c0_U152:Y c0_U152:vdd XNOR2X1
Xc0_U153 c0_U153:A c0_U153:B c0_U153:gnd c0_U153:Y c0_U153:vdd XOR2X1
Xc0_U154 c0_U154:A c0_U154:B c0_U154:gnd c0_U154:Y c0_U154:vdd XNOR2X1
Xc0_U155 c0_U155:A c0_U155:B c0_U155:gnd c0_U155:Y c0_U155:vdd XOR2X1
Xc0_U156 c0_U156:A c0_U156:B c0_U156:gnd c0_U156:Y c0_U156:vdd XNOR2X1
Xc0_U157 c0_U157:A c0_U157:B c0_U157:gnd c0_U157:Y c0_U157:vdd XOR2X1
Xc0_U158 c0_U158:A c0_U158:B c0_U158:gnd c0_U158:Y c0_U158:vdd XNOR2X1
Xc0_U159 c0_U159:A c0_U159:B c0_U159:gnd c0_U159:Y c0_U159:vdd NAND2X1
Xc0_U160 c0_U160:A c0_U160:B c0_U160:gnd c0_U160:Y c0_U160:vdd XOR2X1
Xc0_U161 c0_U161:A c0_U161:B c0_U161:gnd c0_U161:Y c0_U161:vdd XOR2X1
Xc0_U162 c0_U162:A c0_U162:B c0_U162:gnd c0_U162:Y c0_U162:vdd XOR2X1
Xc0_U163 c0_U163:A c0_U163:B c0_U163:gnd c0_U163:Y c0_U163:vdd XOR2X1
Xc0_U164 c0_U164:A c0_U164:B c0_U164:gnd c0_U164:Y c0_U164:vdd XOR2X1
Xc0_U165 c0_U165:A c0_U165:B c0_U165:gnd c0_U165:Y c0_U165:vdd XNOR2X1
Xc0_U166 c0_U166:A c0_U166:B c0_U166:gnd c0_U166:Y c0_U166:vdd XOR2X1
Xc0_U167 c0_U167:A c0_U167:B c0_U167:gnd c0_U167:Y c0_U167:vdd XNOR2X1
Xc0_U168 c0_U168:A c0_U168:B c0_U168:gnd c0_U168:Y c0_U168:vdd XOR2X1
Xc0_U169 c0_U169:A c0_U169:B c0_U169:gnd c0_U169:Y c0_U169:vdd XNOR2X1
Xc0_U170 c0_U170:A c0_U170:B c0_U170:gnd c0_U170:Y c0_U170:vdd XOR2X1
Xc0_U171 c0_U171:A c0_U171:B c0_U171:gnd c0_U171:Y c0_U171:vdd XOR2X1
Xc0_U172 c0_U172:A c0_U172:B c0_U172:gnd c0_U172:Y c0_U172:vdd NAND2X1
Xc0_U173 c0_U173:A c0_U173:B c0_U173:gnd c0_U173:Y c0_U173:vdd XOR2X1
Xc0_U174 c0_U174:A c0_U174:B c0_U174:gnd c0_U174:Y c0_U174:vdd XOR2X1
Xc0_U175 c0_U175:A c0_U175:B c0_U175:gnd c0_U175:Y c0_U175:vdd XOR2X1
Xc0_U176 c0_U176:A c0_U176:B c0_U176:gnd c0_U176:Y c0_U176:vdd XOR2X1
Xc0_U177 c0_U177:A c0_U177:B c0_U177:gnd c0_U177:Y c0_U177:vdd XOR2X1
Xc0_U178 c0_U178:A c0_U178:B c0_U178:gnd c0_U178:Y c0_U178:vdd XNOR2X1
Xc0_U179 c0_U179:A c0_U179:B c0_U179:gnd c0_U179:Y c0_U179:vdd XOR2X1
Xc0_U180 c0_U180:A c0_U180:B c0_U180:gnd c0_U180:Y c0_U180:vdd XOR2X1
Xc0_U181 c0_U181:A c0_U181:B c0_U181:gnd c0_U181:Y c0_U181:vdd XOR2X1
Xc0_U182 c0_U182:A c0_U182:B c0_U182:gnd c0_U182:Y c0_U182:vdd XNOR2X1
Xc0_U183 c0_U183:A c0_U183:B c0_U183:gnd c0_U183:Y c0_U183:vdd XOR2X1
Xc0_U184 c0_U184:A c0_U184:B c0_U184:gnd c0_U184:Y c0_U184:vdd XNOR2X1
Xc0_U185 c0_U185:A c0_U185:B c0_U185:gnd c0_U185:Y c0_U185:vdd NAND2X1
XiDFF_1_q_reg iDFF_1_q_reg:Q iDFF_1_q_reg:CLK iDFF_1_q_reg:D iDFF_1_q_reg:gnd
+  iDFF_1_q_reg:vdd DFFPOSX1
XiDFF_2_q_reg iDFF_2_q_reg:Q iDFF_2_q_reg:CLK iDFF_2_q_reg:D iDFF_2_q_reg:gnd
+  iDFF_2_q_reg:vdd DFFPOSX1
XiDFF_3_q_reg iDFF_3_q_reg:Q iDFF_3_q_reg:CLK iDFF_3_q_reg:D iDFF_3_q_reg:gnd
+  iDFF_3_q_reg:vdd DFFPOSX1
XiDFF_4_q_reg iDFF_4_q_reg:Q iDFF_4_q_reg:CLK iDFF_4_q_reg:D iDFF_4_q_reg:gnd
+  iDFF_4_q_reg:vdd DFFPOSX1
XiDFF_5_q_reg iDFF_5_q_reg:Q iDFF_5_q_reg:CLK iDFF_5_q_reg:D iDFF_5_q_reg:gnd
+  iDFF_5_q_reg:vdd DFFPOSX1
XiDFF_6_q_reg iDFF_6_q_reg:Q iDFF_6_q_reg:CLK iDFF_6_q_reg:D iDFF_6_q_reg:gnd
+  iDFF_6_q_reg:vdd DFFPOSX1
XiDFF_7_q_reg iDFF_7_q_reg:Q iDFF_7_q_reg:CLK iDFF_7_q_reg:D iDFF_7_q_reg:gnd
+  iDFF_7_q_reg:vdd DFFPOSX1
XiDFF_8_q_reg iDFF_8_q_reg:Q iDFF_8_q_reg:CLK iDFF_8_q_reg:D iDFF_8_q_reg:gnd
+  iDFF_8_q_reg:vdd DFFPOSX1
XiDFF_9_q_reg iDFF_9_q_reg:Q iDFF_9_q_reg:CLK iDFF_9_q_reg:D iDFF_9_q_reg:gnd
+  iDFF_9_q_reg:vdd DFFPOSX1
XiDFF_10_q_reg iDFF_10_q_reg:Q iDFF_10_q_reg:CLK iDFF_10_q_reg:D
+  iDFF_10_q_reg:gnd iDFF_10_q_reg:vdd DFFPOSX1
XiDFF_11_q_reg iDFF_11_q_reg:Q iDFF_11_q_reg:CLK iDFF_11_q_reg:D
+  iDFF_11_q_reg:gnd iDFF_11_q_reg:vdd DFFPOSX1
XiDFF_12_q_reg iDFF_12_q_reg:Q iDFF_12_q_reg:CLK iDFF_12_q_reg:D
+  iDFF_12_q_reg:gnd iDFF_12_q_reg:vdd DFFPOSX1
XiDFF_13_q_reg iDFF_13_q_reg:Q iDFF_13_q_reg:CLK iDFF_13_q_reg:D
+  iDFF_13_q_reg:gnd iDFF_13_q_reg:vdd DFFPOSX1
XiDFF_14_q_reg iDFF_14_q_reg:Q iDFF_14_q_reg:CLK iDFF_14_q_reg:D
+  iDFF_14_q_reg:gnd iDFF_14_q_reg:vdd DFFPOSX1
XiDFF_15_q_reg iDFF_15_q_reg:Q iDFF_15_q_reg:CLK iDFF_15_q_reg:D
+  iDFF_15_q_reg:gnd iDFF_15_q_reg:vdd DFFPOSX1
XiDFF_16_q_reg iDFF_16_q_reg:Q iDFF_16_q_reg:CLK iDFF_16_q_reg:D
+  iDFF_16_q_reg:gnd iDFF_16_q_reg:vdd DFFPOSX1
XiDFF_17_q_reg iDFF_17_q_reg:Q iDFF_17_q_reg:CLK iDFF_17_q_reg:D
+  iDFF_17_q_reg:gnd iDFF_17_q_reg:vdd DFFPOSX1
XiDFF_18_q_reg iDFF_18_q_reg:Q iDFF_18_q_reg:CLK iDFF_18_q_reg:D
+  iDFF_18_q_reg:gnd iDFF_18_q_reg:vdd DFFPOSX1
XiDFF_19_q_reg iDFF_19_q_reg:Q iDFF_19_q_reg:CLK iDFF_19_q_reg:D
+  iDFF_19_q_reg:gnd iDFF_19_q_reg:vdd DFFPOSX1
XiDFF_20_q_reg iDFF_20_q_reg:Q iDFF_20_q_reg:CLK iDFF_20_q_reg:D
+  iDFF_20_q_reg:gnd iDFF_20_q_reg:vdd DFFPOSX1
XiDFF_21_q_reg iDFF_21_q_reg:Q iDFF_21_q_reg:CLK iDFF_21_q_reg:D
+  iDFF_21_q_reg:gnd iDFF_21_q_reg:vdd DFFPOSX1
XiDFF_22_q_reg iDFF_22_q_reg:Q iDFF_22_q_reg:CLK iDFF_22_q_reg:D
+  iDFF_22_q_reg:gnd iDFF_22_q_reg:vdd DFFPOSX1
XiDFF_23_q_reg iDFF_23_q_reg:Q iDFF_23_q_reg:CLK iDFF_23_q_reg:D
+  iDFF_23_q_reg:gnd iDFF_23_q_reg:vdd DFFPOSX1
XiDFF_24_q_reg iDFF_24_q_reg:Q iDFF_24_q_reg:CLK iDFF_24_q_reg:D
+  iDFF_24_q_reg:gnd iDFF_24_q_reg:vdd DFFPOSX1
XiDFF_25_q_reg iDFF_25_q_reg:Q iDFF_25_q_reg:CLK iDFF_25_q_reg:D
+  iDFF_25_q_reg:gnd iDFF_25_q_reg:vdd DFFPOSX1
XiDFF_26_q_reg iDFF_26_q_reg:Q iDFF_26_q_reg:CLK iDFF_26_q_reg:D
+  iDFF_26_q_reg:gnd iDFF_26_q_reg:vdd DFFPOSX1
XiDFF_27_q_reg iDFF_27_q_reg:Q iDFF_27_q_reg:CLK iDFF_27_q_reg:D
+  iDFF_27_q_reg:gnd iDFF_27_q_reg:vdd DFFPOSX1
XiDFF_28_q_reg iDFF_28_q_reg:Q iDFF_28_q_reg:CLK iDFF_28_q_reg:D
+  iDFF_28_q_reg:gnd iDFF_28_q_reg:vdd DFFPOSX1
XiDFF_29_q_reg iDFF_29_q_reg:Q iDFF_29_q_reg:CLK iDFF_29_q_reg:D
+  iDFF_29_q_reg:gnd iDFF_29_q_reg:vdd DFFPOSX1
XiDFF_30_q_reg iDFF_30_q_reg:Q iDFF_30_q_reg:CLK iDFF_30_q_reg:D
+  iDFF_30_q_reg:gnd iDFF_30_q_reg:vdd DFFPOSX1
XiDFF_31_q_reg iDFF_31_q_reg:Q iDFF_31_q_reg:CLK iDFF_31_q_reg:D
+  iDFF_31_q_reg:gnd iDFF_31_q_reg:vdd DFFPOSX1
XiDFF_32_q_reg iDFF_32_q_reg:Q iDFF_32_q_reg:CLK iDFF_32_q_reg:D
+  iDFF_32_q_reg:gnd iDFF_32_q_reg:vdd DFFPOSX1
XiDFF_33_q_reg iDFF_33_q_reg:Q iDFF_33_q_reg:CLK iDFF_33_q_reg:D
+  iDFF_33_q_reg:gnd iDFF_33_q_reg:vdd DFFPOSX1
XiDFF_34_q_reg iDFF_34_q_reg:Q iDFF_34_q_reg:CLK iDFF_34_q_reg:D
+  iDFF_34_q_reg:gnd iDFF_34_q_reg:vdd DFFPOSX1
XiDFF_35_q_reg iDFF_35_q_reg:Q iDFF_35_q_reg:CLK iDFF_35_q_reg:D
+  iDFF_35_q_reg:gnd iDFF_35_q_reg:vdd DFFPOSX1
XiDFF_36_q_reg iDFF_36_q_reg:Q iDFF_36_q_reg:CLK iDFF_36_q_reg:D
+  iDFF_36_q_reg:gnd iDFF_36_q_reg:vdd DFFPOSX1
XiDFF_37_q_reg iDFF_37_q_reg:Q iDFF_37_q_reg:CLK iDFF_37_q_reg:D
+  iDFF_37_q_reg:gnd iDFF_37_q_reg:vdd DFFPOSX1
XiDFF_38_q_reg iDFF_38_q_reg:Q iDFF_38_q_reg:CLK iDFF_38_q_reg:D
+  iDFF_38_q_reg:gnd iDFF_38_q_reg:vdd DFFPOSX1
XiDFF_39_q_reg iDFF_39_q_reg:Q iDFF_39_q_reg:CLK iDFF_39_q_reg:D
+  iDFF_39_q_reg:gnd iDFF_39_q_reg:vdd DFFPOSX1
XiDFF_40_q_reg iDFF_40_q_reg:Q iDFF_40_q_reg:CLK iDFF_40_q_reg:D
+  iDFF_40_q_reg:gnd iDFF_40_q_reg:vdd DFFPOSX1
XiDFF_41_q_reg iDFF_41_q_reg:Q iDFF_41_q_reg:CLK iDFF_41_q_reg:D
+  iDFF_41_q_reg:gnd iDFF_41_q_reg:vdd DFFPOSX1
XDFF_1_q_reg DFF_1_q_reg:Q DFF_1_q_reg:CLK DFF_1_q_reg:D DFF_1_q_reg:gnd
+  DFF_1_q_reg:vdd DFFPOSX1
XDFF_2_q_reg DFF_2_q_reg:Q DFF_2_q_reg:CLK DFF_2_q_reg:D DFF_2_q_reg:gnd
+  DFF_2_q_reg:vdd DFFPOSX1
XDFF_3_q_reg DFF_3_q_reg:Q DFF_3_q_reg:CLK DFF_3_q_reg:D DFF_3_q_reg:gnd
+  DFF_3_q_reg:vdd DFFPOSX1
XDFF_4_q_reg DFF_4_q_reg:Q DFF_4_q_reg:CLK DFF_4_q_reg:D DFF_4_q_reg:gnd
+  DFF_4_q_reg:vdd DFFPOSX1
XDFF_5_q_reg DFF_5_q_reg:Q DFF_5_q_reg:CLK DFF_5_q_reg:D DFF_5_q_reg:gnd
+  DFF_5_q_reg:vdd DFFPOSX1
XDFF_6_q_reg DFF_6_q_reg:Q DFF_6_q_reg:CLK DFF_6_q_reg:D DFF_6_q_reg:gnd
+  DFF_6_q_reg:vdd DFFPOSX1
XDFF_7_q_reg DFF_7_q_reg:Q DFF_7_q_reg:CLK DFF_7_q_reg:D DFF_7_q_reg:gnd
+  DFF_7_q_reg:vdd DFFPOSX1
XDFF_8_q_reg DFF_8_q_reg:Q DFF_8_q_reg:CLK DFF_8_q_reg:D DFF_8_q_reg:gnd
+  DFF_8_q_reg:vdd DFFPOSX1
XDFF_9_q_reg DFF_9_q_reg:Q DFF_9_q_reg:CLK DFF_9_q_reg:D DFF_9_q_reg:gnd
+  DFF_9_q_reg:vdd DFFPOSX1
XDFF_10_q_reg DFF_10_q_reg:Q DFF_10_q_reg:CLK DFF_10_q_reg:D DFF_10_q_reg:gnd
+  DFF_10_q_reg:vdd DFFPOSX1
XDFF_11_q_reg DFF_11_q_reg:Q DFF_11_q_reg:CLK DFF_11_q_reg:D DFF_11_q_reg:gnd
+  DFF_11_q_reg:vdd DFFPOSX1
XDFF_12_q_reg DFF_12_q_reg:Q DFF_12_q_reg:CLK DFF_12_q_reg:D DFF_12_q_reg:gnd
+  DFF_12_q_reg:vdd DFFPOSX1
XDFF_13_q_reg DFF_13_q_reg:Q DFF_13_q_reg:CLK DFF_13_q_reg:D DFF_13_q_reg:gnd
+  DFF_13_q_reg:vdd DFFPOSX1
XDFF_14_q_reg DFF_14_q_reg:Q DFF_14_q_reg:CLK DFF_14_q_reg:D DFF_14_q_reg:gnd
+  DFF_14_q_reg:vdd DFFPOSX1
XDFF_15_q_reg DFF_15_q_reg:Q DFF_15_q_reg:CLK DFF_15_q_reg:D DFF_15_q_reg:gnd
+  DFF_15_q_reg:vdd DFFPOSX1
XDFF_16_q_reg DFF_16_q_reg:Q DFF_16_q_reg:CLK DFF_16_q_reg:D DFF_16_q_reg:gnd
+  DFF_16_q_reg:vdd DFFPOSX1
XDFF_17_q_reg DFF_17_q_reg:Q DFF_17_q_reg:CLK DFF_17_q_reg:D DFF_17_q_reg:gnd
+  DFF_17_q_reg:vdd DFFPOSX1
XDFF_18_q_reg DFF_18_q_reg:Q DFF_18_q_reg:CLK DFF_18_q_reg:D DFF_18_q_reg:gnd
+  DFF_18_q_reg:vdd DFFPOSX1
XDFF_19_q_reg DFF_19_q_reg:Q DFF_19_q_reg:CLK DFF_19_q_reg:D DFF_19_q_reg:gnd
+  DFF_19_q_reg:vdd DFFPOSX1
XDFF_20_q_reg DFF_20_q_reg:Q DFF_20_q_reg:CLK DFF_20_q_reg:D DFF_20_q_reg:gnd
+  DFF_20_q_reg:vdd DFFPOSX1
XDFF_21_q_reg DFF_21_q_reg:Q DFF_21_q_reg:CLK DFF_21_q_reg:D DFF_21_q_reg:gnd
+  DFF_21_q_reg:vdd DFFPOSX1
XDFF_22_q_reg DFF_22_q_reg:Q DFF_22_q_reg:CLK DFF_22_q_reg:D DFF_22_q_reg:gnd
+  DFF_22_q_reg:vdd DFFPOSX1
XDFF_23_q_reg DFF_23_q_reg:Q DFF_23_q_reg:CLK DFF_23_q_reg:D DFF_23_q_reg:gnd
+  DFF_23_q_reg:vdd DFFPOSX1
XDFF_24_q_reg DFF_24_q_reg:Q DFF_24_q_reg:CLK DFF_24_q_reg:D DFF_24_q_reg:gnd
+  DFF_24_q_reg:vdd DFFPOSX1
XDFF_25_q_reg DFF_25_q_reg:Q DFF_25_q_reg:CLK DFF_25_q_reg:D DFF_25_q_reg:gnd
+  DFF_25_q_reg:vdd DFFPOSX1
XDFF_26_q_reg DFF_26_q_reg:Q DFF_26_q_reg:CLK DFF_26_q_reg:D DFF_26_q_reg:gnd
+  DFF_26_q_reg:vdd DFFPOSX1
XDFF_27_q_reg DFF_27_q_reg:Q DFF_27_q_reg:CLK DFF_27_q_reg:D DFF_27_q_reg:gnd
+  DFF_27_q_reg:vdd DFFPOSX1
XDFF_28_q_reg DFF_28_q_reg:Q DFF_28_q_reg:CLK DFF_28_q_reg:D DFF_28_q_reg:gnd
+  DFF_28_q_reg:vdd DFFPOSX1
XDFF_29_q_reg DFF_29_q_reg:Q DFF_29_q_reg:CLK DFF_29_q_reg:D DFF_29_q_reg:gnd
+  DFF_29_q_reg:vdd DFFPOSX1
XDFF_30_q_reg DFF_30_q_reg:Q DFF_30_q_reg:CLK DFF_30_q_reg:D DFF_30_q_reg:gnd
+  DFF_30_q_reg:vdd DFFPOSX1
XDFF_31_q_reg DFF_31_q_reg:Q DFF_31_q_reg:CLK DFF_31_q_reg:D DFF_31_q_reg:gnd
+  DFF_31_q_reg:vdd DFFPOSX1
XDFF_32_q_reg DFF_32_q_reg:Q DFF_32_q_reg:CLK DFF_32_q_reg:D DFF_32_q_reg:gnd
+  DFF_32_q_reg:vdd DFFPOSX1
XoDFF_1_q_reg oDFF_1_q_reg:Q oDFF_1_q_reg:CLK oDFF_1_q_reg:D oDFF_1_q_reg:gnd
+  oDFF_1_q_reg:vdd DFFPOSX1
XoDFF_2_q_reg oDFF_2_q_reg:Q oDFF_2_q_reg:CLK oDFF_2_q_reg:D oDFF_2_q_reg:gnd
+  oDFF_2_q_reg:vdd DFFPOSX1
XoDFF_3_q_reg oDFF_3_q_reg:Q oDFF_3_q_reg:CLK oDFF_3_q_reg:D oDFF_3_q_reg:gnd
+  oDFF_3_q_reg:vdd DFFPOSX1
XoDFF_4_q_reg oDFF_4_q_reg:Q oDFF_4_q_reg:CLK oDFF_4_q_reg:D oDFF_4_q_reg:gnd
+  oDFF_4_q_reg:vdd DFFPOSX1
XoDFF_5_q_reg oDFF_5_q_reg:Q oDFF_5_q_reg:CLK oDFF_5_q_reg:D oDFF_5_q_reg:gnd
+  oDFF_5_q_reg:vdd DFFPOSX1
XoDFF_6_q_reg oDFF_6_q_reg:Q oDFF_6_q_reg:CLK oDFF_6_q_reg:D oDFF_6_q_reg:gnd
+  oDFF_6_q_reg:vdd DFFPOSX1
XoDFF_7_q_reg oDFF_7_q_reg:Q oDFF_7_q_reg:CLK oDFF_7_q_reg:D oDFF_7_q_reg:gnd
+  oDFF_7_q_reg:vdd DFFPOSX1
XoDFF_8_q_reg oDFF_8_q_reg:Q oDFF_8_q_reg:CLK oDFF_8_q_reg:D oDFF_8_q_reg:gnd
+  oDFF_8_q_reg:vdd DFFPOSX1
XoDFF_9_q_reg oDFF_9_q_reg:Q oDFF_9_q_reg:CLK oDFF_9_q_reg:D oDFF_9_q_reg:gnd
+  oDFF_9_q_reg:vdd DFFPOSX1
XoDFF_10_q_reg oDFF_10_q_reg:Q oDFF_10_q_reg:CLK oDFF_10_q_reg:D
+  oDFF_10_q_reg:gnd oDFF_10_q_reg:vdd DFFPOSX1
XoDFF_11_q_reg oDFF_11_q_reg:Q oDFF_11_q_reg:CLK oDFF_11_q_reg:D
+  oDFF_11_q_reg:gnd oDFF_11_q_reg:vdd DFFPOSX1
XoDFF_12_q_reg oDFF_12_q_reg:Q oDFF_12_q_reg:CLK oDFF_12_q_reg:D
+  oDFF_12_q_reg:gnd oDFF_12_q_reg:vdd DFFPOSX1
XoDFF_13_q_reg oDFF_13_q_reg:Q oDFF_13_q_reg:CLK oDFF_13_q_reg:D
+  oDFF_13_q_reg:gnd oDFF_13_q_reg:vdd DFFPOSX1
XoDFF_14_q_reg oDFF_14_q_reg:Q oDFF_14_q_reg:CLK oDFF_14_q_reg:D
+  oDFF_14_q_reg:gnd oDFF_14_q_reg:vdd DFFPOSX1
XoDFF_15_q_reg oDFF_15_q_reg:Q oDFF_15_q_reg:CLK oDFF_15_q_reg:D
+  oDFF_15_q_reg:gnd oDFF_15_q_reg:vdd DFFPOSX1
XoDFF_16_q_reg oDFF_16_q_reg:Q oDFF_16_q_reg:CLK oDFF_16_q_reg:D
+  oDFF_16_q_reg:gnd oDFF_16_q_reg:vdd DFFPOSX1
XoDFF_17_q_reg oDFF_17_q_reg:Q oDFF_17_q_reg:CLK oDFF_17_q_reg:D
+  oDFF_17_q_reg:gnd oDFF_17_q_reg:vdd DFFPOSX1
XoDFF_18_q_reg oDFF_18_q_reg:Q oDFF_18_q_reg:CLK oDFF_18_q_reg:D
+  oDFF_18_q_reg:gnd oDFF_18_q_reg:vdd DFFPOSX1
XoDFF_19_q_reg oDFF_19_q_reg:Q oDFF_19_q_reg:CLK oDFF_19_q_reg:D
+  oDFF_19_q_reg:gnd oDFF_19_q_reg:vdd DFFPOSX1
XoDFF_20_q_reg oDFF_20_q_reg:Q oDFF_20_q_reg:CLK oDFF_20_q_reg:D
+  oDFF_20_q_reg:gnd oDFF_20_q_reg:vdd DFFPOSX1
XoDFF_21_q_reg oDFF_21_q_reg:Q oDFF_21_q_reg:CLK oDFF_21_q_reg:D
+  oDFF_21_q_reg:gnd oDFF_21_q_reg:vdd DFFPOSX1
XoDFF_22_q_reg oDFF_22_q_reg:Q oDFF_22_q_reg:CLK oDFF_22_q_reg:D
+  oDFF_22_q_reg:gnd oDFF_22_q_reg:vdd DFFPOSX1
XoDFF_23_q_reg oDFF_23_q_reg:Q oDFF_23_q_reg:CLK oDFF_23_q_reg:D
+  oDFF_23_q_reg:gnd oDFF_23_q_reg:vdd DFFPOSX1
XoDFF_24_q_reg oDFF_24_q_reg:Q oDFF_24_q_reg:CLK oDFF_24_q_reg:D
+  oDFF_24_q_reg:gnd oDFF_24_q_reg:vdd DFFPOSX1
XoDFF_25_q_reg oDFF_25_q_reg:Q oDFF_25_q_reg:CLK oDFF_25_q_reg:D
+  oDFF_25_q_reg:gnd oDFF_25_q_reg:vdd DFFPOSX1
XoDFF_26_q_reg oDFF_26_q_reg:Q oDFF_26_q_reg:CLK oDFF_26_q_reg:D
+  oDFF_26_q_reg:gnd oDFF_26_q_reg:vdd DFFPOSX1
XoDFF_27_q_reg oDFF_27_q_reg:Q oDFF_27_q_reg:CLK oDFF_27_q_reg:D
+  oDFF_27_q_reg:gnd oDFF_27_q_reg:vdd DFFPOSX1
XoDFF_28_q_reg oDFF_28_q_reg:Q oDFF_28_q_reg:CLK oDFF_28_q_reg:D
+  oDFF_28_q_reg:gnd oDFF_28_q_reg:vdd DFFPOSX1
XoDFF_29_q_reg oDFF_29_q_reg:Q oDFF_29_q_reg:CLK oDFF_29_q_reg:D
+  oDFF_29_q_reg:gnd oDFF_29_q_reg:vdd DFFPOSX1
XoDFF_30_q_reg oDFF_30_q_reg:Q oDFF_30_q_reg:CLK oDFF_30_q_reg:D
+  oDFF_30_q_reg:gnd oDFF_30_q_reg:vdd DFFPOSX1
XoDFF_31_q_reg oDFF_31_q_reg:Q oDFF_31_q_reg:CLK oDFF_31_q_reg:D
+  oDFF_31_q_reg:gnd oDFF_31_q_reg:vdd DFFPOSX1
XoDFF_32_q_reg oDFF_32_q_reg:Q oDFF_32_q_reg:CLK oDFF_32_q_reg:D
+  oDFF_32_q_reg:gnd oDFF_32_q_reg:vdd DFFPOSX1
.ENDS


******Simulation parameters*****

****Param definitions***
.param clk_period= '(1/100)*(0.000001)' 
+half_clk_period= '(clk_period/2)'
+double_clk_period= '(clk_period*2)'

.param fall_from_value=6e-08
+ fall_to_value=6.2e-08

.param init_delay = half_clk_period
+ rise_time= 50p
+ fall_time= 50p

.param change_time='(half_clk_period/3)'
.param k_minus_4='(half_clk_period/3)'
.param k_minus_3='k_minus_4 + clk_period'
.param k_minus_3rise='k_minus_3 + 100ps'
.param k_minus_2='k_minus_3 + clk_period'
.param k_minus_2rise='k_minus_2 + 100ps'
.param k_minus_1='k_minus_2 + clk_period'
.param k_minus_1rise='k_minus_1 + 100ps'
.param k_cycle = 'k_minus_1 + clk_period'
.param k_cycle_rise = 'k_cycle + 100ps'
.param k_plus1= '(k_cycle + half_clk_period )'
.param k_plus1_rise = '(k_plus1 + 100ps)'
.param current_magnitude = 2.2mA
+rise_delay= ##glitch_location##s
+fall_delay= 'rise_delay+5p'
+rise_time_constant = 1ps
+fall_time_constant=130ps

.GLOBAL vdd VDD

Vvdd vdd 0 1.8
VCk  clk   0  PULSE(0 1.8 init_delay rise_time fall_time half_clk_period clk_period)



******Instantiating the subckt*****

Xc499_clk_opFF
+       clk N1 N5 N9 N13 N17 N21 N25 N29 N33 N37 N41 N45 N49 N53 N57 N61 N65 N69
+       N73 N77 N81 N85 N89 N93 N97 N101 N105 N109 N113 N117 N121 N125 N129 N130
+       N131 N132 N133 N134 N135 N136 N137 Qout_N724 Qout_N725 Qout_N726
+       Qout_N727 Qout_N728 Qout_N729 Qout_N730 Qout_N731 Qout_N732 Qout_N733
+       Qout_N734 Qout_N735 Qout_N736 Qout_N737 Qout_N738 Qout_N739 Qout_N740
+       Qout_N741 Qout_N742 Qout_N743 Qout_N744 Qout_N745 Qout_N746 Qout_N747
+       Qout_N748 Qout_N749 Qout_N750 Qout_N751 Qout_N752 Qout_N753 Qout_N754
+       Qout_N755 c499_clk_opFF

******Done instantiating the subckt*****


V1 N1 0 PWL( 0 ##N1_reference_minus4##  k_minus_3 ##N1_reference_minus4## k_minus_3rise ##N1_reference_minus3## k_minus_2 ##N1_reference_minus3## k_minus_2rise ##N1_reference_minus2## k_minus_1 ##N1_reference_minus2## k_minus_1rise ##N1_reference_minus1## k_cycle ##N1_reference_minus1## k_cycle_rise ##N1_reference_1## k_plus1 ##N1_reference_1## k_plus1_rise ##N1_reference_2## 6.5e-08 ##N1_reference_2##)


V2 N5 0 PWL( 0 ##N5_reference_minus4##  k_minus_3 ##N5_reference_minus4## k_minus_3rise ##N5_reference_minus3## k_minus_2 ##N5_reference_minus3## k_minus_2rise ##N5_reference_minus2## k_minus_1 ##N5_reference_minus2## k_minus_1rise ##N5_reference_minus1## k_cycle ##N5_reference_minus1## k_cycle_rise ##N5_reference_1## k_plus1 ##N5_reference_1## k_plus1_rise ##N5_reference_2## 6.5e-08 ##N5_reference_2##)


V3 N9 0 PWL( 0 ##N9_reference_minus4##  k_minus_3 ##N9_reference_minus4## k_minus_3rise ##N9_reference_minus3## k_minus_2 ##N9_reference_minus3## k_minus_2rise ##N9_reference_minus2## k_minus_1 ##N9_reference_minus2## k_minus_1rise ##N9_reference_minus1## k_cycle ##N9_reference_minus1## k_cycle_rise ##N9_reference_1## k_plus1 ##N9_reference_1## k_plus1_rise ##N9_reference_2## 6.5e-08 ##N9_reference_2##)


V4 N13 0 PWL( 0 ##N13_reference_minus4##  k_minus_3 ##N13_reference_minus4## k_minus_3rise ##N13_reference_minus3## k_minus_2 ##N13_reference_minus3## k_minus_2rise ##N13_reference_minus2## k_minus_1 ##N13_reference_minus2## k_minus_1rise ##N13_reference_minus1## k_cycle ##N13_reference_minus1## k_cycle_rise ##N13_reference_1## k_plus1 ##N13_reference_1## k_plus1_rise ##N13_reference_2## 6.5e-08 ##N13_reference_2##)


V5 N17 0 PWL( 0 ##N17_reference_minus4##  k_minus_3 ##N17_reference_minus4## k_minus_3rise ##N17_reference_minus3## k_minus_2 ##N17_reference_minus3## k_minus_2rise ##N17_reference_minus2## k_minus_1 ##N17_reference_minus2## k_minus_1rise ##N17_reference_minus1## k_cycle ##N17_reference_minus1## k_cycle_rise ##N17_reference_1## k_plus1 ##N17_reference_1## k_plus1_rise ##N17_reference_2## 6.5e-08 ##N17_reference_2##)


V6 N21 0 PWL( 0 ##N21_reference_minus4##  k_minus_3 ##N21_reference_minus4## k_minus_3rise ##N21_reference_minus3## k_minus_2 ##N21_reference_minus3## k_minus_2rise ##N21_reference_minus2## k_minus_1 ##N21_reference_minus2## k_minus_1rise ##N21_reference_minus1## k_cycle ##N21_reference_minus1## k_cycle_rise ##N21_reference_1## k_plus1 ##N21_reference_1## k_plus1_rise ##N21_reference_2## 6.5e-08 ##N21_reference_2##)


V7 N25 0 PWL( 0 ##N25_reference_minus4##  k_minus_3 ##N25_reference_minus4## k_minus_3rise ##N25_reference_minus3## k_minus_2 ##N25_reference_minus3## k_minus_2rise ##N25_reference_minus2## k_minus_1 ##N25_reference_minus2## k_minus_1rise ##N25_reference_minus1## k_cycle ##N25_reference_minus1## k_cycle_rise ##N25_reference_1## k_plus1 ##N25_reference_1## k_plus1_rise ##N25_reference_2## 6.5e-08 ##N25_reference_2##)


V8 N29 0 PWL( 0 ##N29_reference_minus4##  k_minus_3 ##N29_reference_minus4## k_minus_3rise ##N29_reference_minus3## k_minus_2 ##N29_reference_minus3## k_minus_2rise ##N29_reference_minus2## k_minus_1 ##N29_reference_minus2## k_minus_1rise ##N29_reference_minus1## k_cycle ##N29_reference_minus1## k_cycle_rise ##N29_reference_1## k_plus1 ##N29_reference_1## k_plus1_rise ##N29_reference_2## 6.5e-08 ##N29_reference_2##)


V9 N33 0 PWL( 0 ##N33_reference_minus4##  k_minus_3 ##N33_reference_minus4## k_minus_3rise ##N33_reference_minus3## k_minus_2 ##N33_reference_minus3## k_minus_2rise ##N33_reference_minus2## k_minus_1 ##N33_reference_minus2## k_minus_1rise ##N33_reference_minus1## k_cycle ##N33_reference_minus1## k_cycle_rise ##N33_reference_1## k_plus1 ##N33_reference_1## k_plus1_rise ##N33_reference_2## 6.5e-08 ##N33_reference_2##)


V10 N37 0 PWL( 0 ##N37_reference_minus4##  k_minus_3 ##N37_reference_minus4## k_minus_3rise ##N37_reference_minus3## k_minus_2 ##N37_reference_minus3## k_minus_2rise ##N37_reference_minus2## k_minus_1 ##N37_reference_minus2## k_minus_1rise ##N37_reference_minus1## k_cycle ##N37_reference_minus1## k_cycle_rise ##N37_reference_1## k_plus1 ##N37_reference_1## k_plus1_rise ##N37_reference_2## 6.5e-08 ##N37_reference_2##)


V11 N41 0 PWL( 0 ##N41_reference_minus4##  k_minus_3 ##N41_reference_minus4## k_minus_3rise ##N41_reference_minus3## k_minus_2 ##N41_reference_minus3## k_minus_2rise ##N41_reference_minus2## k_minus_1 ##N41_reference_minus2## k_minus_1rise ##N41_reference_minus1## k_cycle ##N41_reference_minus1## k_cycle_rise ##N41_reference_1## k_plus1 ##N41_reference_1## k_plus1_rise ##N41_reference_2## 6.5e-08 ##N41_reference_2##)


V12 N45 0 PWL( 0 ##N45_reference_minus4##  k_minus_3 ##N45_reference_minus4## k_minus_3rise ##N45_reference_minus3## k_minus_2 ##N45_reference_minus3## k_minus_2rise ##N45_reference_minus2## k_minus_1 ##N45_reference_minus2## k_minus_1rise ##N45_reference_minus1## k_cycle ##N45_reference_minus1## k_cycle_rise ##N45_reference_1## k_plus1 ##N45_reference_1## k_plus1_rise ##N45_reference_2## 6.5e-08 ##N45_reference_2##)


V13 N49 0 PWL( 0 ##N49_reference_minus4##  k_minus_3 ##N49_reference_minus4## k_minus_3rise ##N49_reference_minus3## k_minus_2 ##N49_reference_minus3## k_minus_2rise ##N49_reference_minus2## k_minus_1 ##N49_reference_minus2## k_minus_1rise ##N49_reference_minus1## k_cycle ##N49_reference_minus1## k_cycle_rise ##N49_reference_1## k_plus1 ##N49_reference_1## k_plus1_rise ##N49_reference_2## 6.5e-08 ##N49_reference_2##)


V14 N53 0 PWL( 0 ##N53_reference_minus4##  k_minus_3 ##N53_reference_minus4## k_minus_3rise ##N53_reference_minus3## k_minus_2 ##N53_reference_minus3## k_minus_2rise ##N53_reference_minus2## k_minus_1 ##N53_reference_minus2## k_minus_1rise ##N53_reference_minus1## k_cycle ##N53_reference_minus1## k_cycle_rise ##N53_reference_1## k_plus1 ##N53_reference_1## k_plus1_rise ##N53_reference_2## 6.5e-08 ##N53_reference_2##)


V15 N57 0 PWL( 0 ##N57_reference_minus4##  k_minus_3 ##N57_reference_minus4## k_minus_3rise ##N57_reference_minus3## k_minus_2 ##N57_reference_minus3## k_minus_2rise ##N57_reference_minus2## k_minus_1 ##N57_reference_minus2## k_minus_1rise ##N57_reference_minus1## k_cycle ##N57_reference_minus1## k_cycle_rise ##N57_reference_1## k_plus1 ##N57_reference_1## k_plus1_rise ##N57_reference_2## 6.5e-08 ##N57_reference_2##)


V16 N61 0 PWL( 0 ##N61_reference_minus4##  k_minus_3 ##N61_reference_minus4## k_minus_3rise ##N61_reference_minus3## k_minus_2 ##N61_reference_minus3## k_minus_2rise ##N61_reference_minus2## k_minus_1 ##N61_reference_minus2## k_minus_1rise ##N61_reference_minus1## k_cycle ##N61_reference_minus1## k_cycle_rise ##N61_reference_1## k_plus1 ##N61_reference_1## k_plus1_rise ##N61_reference_2## 6.5e-08 ##N61_reference_2##)


V17 N65 0 PWL( 0 ##N65_reference_minus4##  k_minus_3 ##N65_reference_minus4## k_minus_3rise ##N65_reference_minus3## k_minus_2 ##N65_reference_minus3## k_minus_2rise ##N65_reference_minus2## k_minus_1 ##N65_reference_minus2## k_minus_1rise ##N65_reference_minus1## k_cycle ##N65_reference_minus1## k_cycle_rise ##N65_reference_1## k_plus1 ##N65_reference_1## k_plus1_rise ##N65_reference_2## 6.5e-08 ##N65_reference_2##)


V18 N69 0 PWL( 0 ##N69_reference_minus4##  k_minus_3 ##N69_reference_minus4## k_minus_3rise ##N69_reference_minus3## k_minus_2 ##N69_reference_minus3## k_minus_2rise ##N69_reference_minus2## k_minus_1 ##N69_reference_minus2## k_minus_1rise ##N69_reference_minus1## k_cycle ##N69_reference_minus1## k_cycle_rise ##N69_reference_1## k_plus1 ##N69_reference_1## k_plus1_rise ##N69_reference_2## 6.5e-08 ##N69_reference_2##)


V19 N73 0 PWL( 0 ##N73_reference_minus4##  k_minus_3 ##N73_reference_minus4## k_minus_3rise ##N73_reference_minus3## k_minus_2 ##N73_reference_minus3## k_minus_2rise ##N73_reference_minus2## k_minus_1 ##N73_reference_minus2## k_minus_1rise ##N73_reference_minus1## k_cycle ##N73_reference_minus1## k_cycle_rise ##N73_reference_1## k_plus1 ##N73_reference_1## k_plus1_rise ##N73_reference_2## 6.5e-08 ##N73_reference_2##)


V20 N77 0 PWL( 0 ##N77_reference_minus4##  k_minus_3 ##N77_reference_minus4## k_minus_3rise ##N77_reference_minus3## k_minus_2 ##N77_reference_minus3## k_minus_2rise ##N77_reference_minus2## k_minus_1 ##N77_reference_minus2## k_minus_1rise ##N77_reference_minus1## k_cycle ##N77_reference_minus1## k_cycle_rise ##N77_reference_1## k_plus1 ##N77_reference_1## k_plus1_rise ##N77_reference_2## 6.5e-08 ##N77_reference_2##)


V21 N81 0 PWL( 0 ##N81_reference_minus4##  k_minus_3 ##N81_reference_minus4## k_minus_3rise ##N81_reference_minus3## k_minus_2 ##N81_reference_minus3## k_minus_2rise ##N81_reference_minus2## k_minus_1 ##N81_reference_minus2## k_minus_1rise ##N81_reference_minus1## k_cycle ##N81_reference_minus1## k_cycle_rise ##N81_reference_1## k_plus1 ##N81_reference_1## k_plus1_rise ##N81_reference_2## 6.5e-08 ##N81_reference_2##)


V22 N85 0 PWL( 0 ##N85_reference_minus4##  k_minus_3 ##N85_reference_minus4## k_minus_3rise ##N85_reference_minus3## k_minus_2 ##N85_reference_minus3## k_minus_2rise ##N85_reference_minus2## k_minus_1 ##N85_reference_minus2## k_minus_1rise ##N85_reference_minus1## k_cycle ##N85_reference_minus1## k_cycle_rise ##N85_reference_1## k_plus1 ##N85_reference_1## k_plus1_rise ##N85_reference_2## 6.5e-08 ##N85_reference_2##)


V23 N89 0 PWL( 0 ##N89_reference_minus4##  k_minus_3 ##N89_reference_minus4## k_minus_3rise ##N89_reference_minus3## k_minus_2 ##N89_reference_minus3## k_minus_2rise ##N89_reference_minus2## k_minus_1 ##N89_reference_minus2## k_minus_1rise ##N89_reference_minus1## k_cycle ##N89_reference_minus1## k_cycle_rise ##N89_reference_1## k_plus1 ##N89_reference_1## k_plus1_rise ##N89_reference_2## 6.5e-08 ##N89_reference_2##)


V24 N93 0 PWL( 0 ##N93_reference_minus4##  k_minus_3 ##N93_reference_minus4## k_minus_3rise ##N93_reference_minus3## k_minus_2 ##N93_reference_minus3## k_minus_2rise ##N93_reference_minus2## k_minus_1 ##N93_reference_minus2## k_minus_1rise ##N93_reference_minus1## k_cycle ##N93_reference_minus1## k_cycle_rise ##N93_reference_1## k_plus1 ##N93_reference_1## k_plus1_rise ##N93_reference_2## 6.5e-08 ##N93_reference_2##)


V25 N97 0 PWL( 0 ##N97_reference_minus4##  k_minus_3 ##N97_reference_minus4## k_minus_3rise ##N97_reference_minus3## k_minus_2 ##N97_reference_minus3## k_minus_2rise ##N97_reference_minus2## k_minus_1 ##N97_reference_minus2## k_minus_1rise ##N97_reference_minus1## k_cycle ##N97_reference_minus1## k_cycle_rise ##N97_reference_1## k_plus1 ##N97_reference_1## k_plus1_rise ##N97_reference_2## 6.5e-08 ##N97_reference_2##)


V26 N101 0 PWL( 0 ##N101_reference_minus4##  k_minus_3 ##N101_reference_minus4## k_minus_3rise ##N101_reference_minus3## k_minus_2 ##N101_reference_minus3## k_minus_2rise ##N101_reference_minus2## k_minus_1 ##N101_reference_minus2## k_minus_1rise ##N101_reference_minus1## k_cycle ##N101_reference_minus1## k_cycle_rise ##N101_reference_1## k_plus1 ##N101_reference_1## k_plus1_rise ##N101_reference_2## 6.5e-08 ##N101_reference_2##)


V27 N105 0 PWL( 0 ##N105_reference_minus4##  k_minus_3 ##N105_reference_minus4## k_minus_3rise ##N105_reference_minus3## k_minus_2 ##N105_reference_minus3## k_minus_2rise ##N105_reference_minus2## k_minus_1 ##N105_reference_minus2## k_minus_1rise ##N105_reference_minus1## k_cycle ##N105_reference_minus1## k_cycle_rise ##N105_reference_1## k_plus1 ##N105_reference_1## k_plus1_rise ##N105_reference_2## 6.5e-08 ##N105_reference_2##)


V28 N109 0 PWL( 0 ##N109_reference_minus4##  k_minus_3 ##N109_reference_minus4## k_minus_3rise ##N109_reference_minus3## k_minus_2 ##N109_reference_minus3## k_minus_2rise ##N109_reference_minus2## k_minus_1 ##N109_reference_minus2## k_minus_1rise ##N109_reference_minus1## k_cycle ##N109_reference_minus1## k_cycle_rise ##N109_reference_1## k_plus1 ##N109_reference_1## k_plus1_rise ##N109_reference_2## 6.5e-08 ##N109_reference_2##)


V29 N113 0 PWL( 0 ##N113_reference_minus4##  k_minus_3 ##N113_reference_minus4## k_minus_3rise ##N113_reference_minus3## k_minus_2 ##N113_reference_minus3## k_minus_2rise ##N113_reference_minus2## k_minus_1 ##N113_reference_minus2## k_minus_1rise ##N113_reference_minus1## k_cycle ##N113_reference_minus1## k_cycle_rise ##N113_reference_1## k_plus1 ##N113_reference_1## k_plus1_rise ##N113_reference_2## 6.5e-08 ##N113_reference_2##)


V30 N117 0 PWL( 0 ##N117_reference_minus4##  k_minus_3 ##N117_reference_minus4## k_minus_3rise ##N117_reference_minus3## k_minus_2 ##N117_reference_minus3## k_minus_2rise ##N117_reference_minus2## k_minus_1 ##N117_reference_minus2## k_minus_1rise ##N117_reference_minus1## k_cycle ##N117_reference_minus1## k_cycle_rise ##N117_reference_1## k_plus1 ##N117_reference_1## k_plus1_rise ##N117_reference_2## 6.5e-08 ##N117_reference_2##)


V31 N121 0 PWL( 0 ##N121_reference_minus4##  k_minus_3 ##N121_reference_minus4## k_minus_3rise ##N121_reference_minus3## k_minus_2 ##N121_reference_minus3## k_minus_2rise ##N121_reference_minus2## k_minus_1 ##N121_reference_minus2## k_minus_1rise ##N121_reference_minus1## k_cycle ##N121_reference_minus1## k_cycle_rise ##N121_reference_1## k_plus1 ##N121_reference_1## k_plus1_rise ##N121_reference_2## 6.5e-08 ##N121_reference_2##)


V32 N125 0 PWL( 0 ##N125_reference_minus4##  k_minus_3 ##N125_reference_minus4## k_minus_3rise ##N125_reference_minus3## k_minus_2 ##N125_reference_minus3## k_minus_2rise ##N125_reference_minus2## k_minus_1 ##N125_reference_minus2## k_minus_1rise ##N125_reference_minus1## k_cycle ##N125_reference_minus1## k_cycle_rise ##N125_reference_1## k_plus1 ##N125_reference_1## k_plus1_rise ##N125_reference_2## 6.5e-08 ##N125_reference_2##)


V33 N129 0 PWL( 0 ##N129_reference_minus4##  k_minus_3 ##N129_reference_minus4## k_minus_3rise ##N129_reference_minus3## k_minus_2 ##N129_reference_minus3## k_minus_2rise ##N129_reference_minus2## k_minus_1 ##N129_reference_minus2## k_minus_1rise ##N129_reference_minus1## k_cycle ##N129_reference_minus1## k_cycle_rise ##N129_reference_1## k_plus1 ##N129_reference_1## k_plus1_rise ##N129_reference_2## 6.5e-08 ##N129_reference_2##)


V34 N130 0 PWL( 0 ##N130_reference_minus4##  k_minus_3 ##N130_reference_minus4## k_minus_3rise ##N130_reference_minus3## k_minus_2 ##N130_reference_minus3## k_minus_2rise ##N130_reference_minus2## k_minus_1 ##N130_reference_minus2## k_minus_1rise ##N130_reference_minus1## k_cycle ##N130_reference_minus1## k_cycle_rise ##N130_reference_1## k_plus1 ##N130_reference_1## k_plus1_rise ##N130_reference_2## 6.5e-08 ##N130_reference_2##)


V35 N131 0 PWL( 0 ##N131_reference_minus4##  k_minus_3 ##N131_reference_minus4## k_minus_3rise ##N131_reference_minus3## k_minus_2 ##N131_reference_minus3## k_minus_2rise ##N131_reference_minus2## k_minus_1 ##N131_reference_minus2## k_minus_1rise ##N131_reference_minus1## k_cycle ##N131_reference_minus1## k_cycle_rise ##N131_reference_1## k_plus1 ##N131_reference_1## k_plus1_rise ##N131_reference_2## 6.5e-08 ##N131_reference_2##)


V36 N132 0 PWL( 0 ##N132_reference_minus4##  k_minus_3 ##N132_reference_minus4## k_minus_3rise ##N132_reference_minus3## k_minus_2 ##N132_reference_minus3## k_minus_2rise ##N132_reference_minus2## k_minus_1 ##N132_reference_minus2## k_minus_1rise ##N132_reference_minus1## k_cycle ##N132_reference_minus1## k_cycle_rise ##N132_reference_1## k_plus1 ##N132_reference_1## k_plus1_rise ##N132_reference_2## 6.5e-08 ##N132_reference_2##)


V37 N133 0 PWL( 0 ##N133_reference_minus4##  k_minus_3 ##N133_reference_minus4## k_minus_3rise ##N133_reference_minus3## k_minus_2 ##N133_reference_minus3## k_minus_2rise ##N133_reference_minus2## k_minus_1 ##N133_reference_minus2## k_minus_1rise ##N133_reference_minus1## k_cycle ##N133_reference_minus1## k_cycle_rise ##N133_reference_1## k_plus1 ##N133_reference_1## k_plus1_rise ##N133_reference_2## 6.5e-08 ##N133_reference_2##)


V38 N134 0 PWL( 0 ##N134_reference_minus4##  k_minus_3 ##N134_reference_minus4## k_minus_3rise ##N134_reference_minus3## k_minus_2 ##N134_reference_minus3## k_minus_2rise ##N134_reference_minus2## k_minus_1 ##N134_reference_minus2## k_minus_1rise ##N134_reference_minus1## k_cycle ##N134_reference_minus1## k_cycle_rise ##N134_reference_1## k_plus1 ##N134_reference_1## k_plus1_rise ##N134_reference_2## 6.5e-08 ##N134_reference_2##)


V39 N135 0 PWL( 0 ##N135_reference_minus4##  k_minus_3 ##N135_reference_minus4## k_minus_3rise ##N135_reference_minus3## k_minus_2 ##N135_reference_minus3## k_minus_2rise ##N135_reference_minus2## k_minus_1 ##N135_reference_minus2## k_minus_1rise ##N135_reference_minus1## k_cycle ##N135_reference_minus1## k_cycle_rise ##N135_reference_1## k_plus1 ##N135_reference_1## k_plus1_rise ##N135_reference_2## 6.5e-08 ##N135_reference_2##)


V40 N136 0 PWL( 0 ##N136_reference_minus4##  k_minus_3 ##N136_reference_minus4## k_minus_3rise ##N136_reference_minus3## k_minus_2 ##N136_reference_minus3## k_minus_2rise ##N136_reference_minus2## k_minus_1 ##N136_reference_minus2## k_minus_1rise ##N136_reference_minus1## k_cycle ##N136_reference_minus1## k_cycle_rise ##N136_reference_1## k_plus1 ##N136_reference_1## k_plus1_rise ##N136_reference_2## 6.5e-08 ##N136_reference_2##)


V41 N137 0 PWL( 0 ##N137_reference_minus4##  k_minus_3 ##N137_reference_minus4## k_minus_3rise ##N137_reference_minus3## k_minus_2 ##N137_reference_minus3## k_minus_2rise ##N137_reference_minus2## k_minus_1 ##N137_reference_minus2## k_minus_1rise ##N137_reference_minus1## k_cycle ##N137_reference_minus1## k_cycle_rise ##N137_reference_1## k_plus1 ##N137_reference_1## k_plus1_rise ##N137_reference_2## 6.5e-08 ##N137_reference_2##)

**Initialising input of all FFs- commented this out. Doesnt help.PWL

**Initialising output of all FFs- trying..

*.ic v(Xc499_clk_opFF.iDFF_1:Q)= ##IN_N1_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_2:Q)= ##IN_N5_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_3:Q)= ##IN_N9_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_4:Q)= ##IN_N13_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_5:Q)= ##IN_N17_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_6:Q)= ##IN_N21_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_7:Q)= ##IN_N25_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_8:Q)= ##IN_N29_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_9:Q)= ##IN_N33_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_10:Q)= ##IN_N37_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_11:Q)= ##IN_N41_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_12:Q)= ##IN_N45_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_13:Q)= ##IN_N49_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_14:Q)= ##IN_N53_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_15:Q)= ##IN_N57_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_16:Q)= ##IN_N61_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_17:Q)= ##IN_N65_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_18:Q)= ##IN_N69_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_19:Q)= ##IN_N73_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_20:Q)= ##IN_N77_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_21:Q)= ##IN_N81_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_22:Q)= ##IN_N85_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_23:Q)= ##IN_N89_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_24:Q)= ##IN_N93_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_25:Q)= ##IN_N97_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_26:Q)= ##IN_N101_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_27:Q)= ##IN_N105_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_28:Q)= ##IN_N109_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_29:Q)= ##IN_N113_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_30:Q)= ##IN_N117_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_31:Q)= ##IN_N121_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_32:Q)= ##IN_N125_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_33:Q)= ##IN_N129_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_34:Q)= ##IN_N130_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_35:Q)= ##IN_N131_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_36:Q)= ##IN_N132_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_37:Q)= ##IN_N133_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_38:Q)= ##IN_N134_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_39:Q)= ##IN_N135_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_40:Q)= ##IN_N136_reference_minus5##
*.ic v(Xc499_clk_opFF.iDFF_41:Q)= ##IN_N137_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_1:Q)= ##Q_N724_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_2:Q)= ##Q_N725_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_3:Q)= ##Q_N726_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_4:Q)= ##Q_N727_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_5:Q)= ##Q_N728_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_6:Q)= ##Q_N729_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_7:Q)= ##Q_N730_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_8:Q)= ##Q_N731_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_9:Q)= ##Q_N732_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_10:Q)= ##Q_N733_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_11:Q)= ##Q_N734_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_12:Q)= ##Q_N735_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_13:Q)= ##Q_N736_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_14:Q)= ##Q_N737_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_15:Q)= ##Q_N738_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_16:Q)= ##Q_N739_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_17:Q)= ##Q_N740_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_18:Q)= ##Q_N741_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_19:Q)= ##Q_N742_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_20:Q)= ##Q_N743_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_21:Q)= ##Q_N744_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_22:Q)= ##Q_N745_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_23:Q)= ##Q_N746_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_24:Q)= ##Q_N747_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_25:Q)= ##Q_N748_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_26:Q)= ##Q_N749_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_27:Q)= ##Q_N750_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_28:Q)= ##Q_N751_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_29:Q)= ##Q_N752_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_30:Q)= ##Q_N753_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_31:Q)= ##Q_N754_reference_minus5##
*.ic v(Xc499_clk_opFF.DFF_32:Q)= ##Q_N755_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_1:Q)= ##Qout_N724_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_2:Q)= ##Qout_N725_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_3:Q)= ##Qout_N726_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_4:Q)= ##Qout_N727_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_5:Q)= ##Qout_N728_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_6:Q)= ##Qout_N729_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_7:Q)= ##Qout_N730_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_8:Q)= ##Qout_N731_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_9:Q)= ##Qout_N732_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_10:Q)= ##Qout_N733_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_11:Q)= ##Qout_N734_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_12:Q)= ##Qout_N735_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_13:Q)= ##Qout_N736_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_14:Q)= ##Qout_N737_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_15:Q)= ##Qout_N738_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_16:Q)= ##Qout_N739_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_17:Q)= ##Qout_N740_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_18:Q)= ##Qout_N741_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_19:Q)= ##Qout_N742_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_20:Q)= ##Qout_N743_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_21:Q)= ##Qout_N744_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_22:Q)= ##Qout_N745_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_23:Q)= ##Qout_N746_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_24:Q)= ##Qout_N747_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_25:Q)= ##Qout_N748_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_26:Q)= ##Qout_N749_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_27:Q)= ##Qout_N750_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_28:Q)= ##Qout_N751_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_29:Q)= ##Qout_N752_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_30:Q)= ##Qout_N753_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_31:Q)= ##Qout_N754_reference_minus5##
*.ic v(Xc499_clk_opFF.oDFF_32:Q)= ##Qout_N755_reference_minus5##

**Initialising primary outputs

*.ic v(Qout_N724)= 0
*.ic v(Qout_N725)= 0
*.ic v(Qout_N726)= 0
*.ic v(Qout_N727)= 0
*.ic v(Qout_N728)= 0
*.ic v(Qout_N729)= 0
*.ic v(Qout_N730)= 0
*.ic v(Qout_N731)= 0
*.ic v(Qout_N732)= 0
*.ic v(Qout_N733)= 0
*.ic v(Qout_N734)= 0
*.ic v(Qout_N735)= 0
*.ic v(Qout_N736)= 0
*.ic v(Qout_N737)= 0
*.ic v(Qout_N738)= 0
*.ic v(Qout_N739)= 0
*.ic v(Qout_N740)= 0
*.ic v(Qout_N741)= 0
*.ic v(Qout_N742)= 0
*.ic v(Qout_N743)= 0
*.ic v(Qout_N744)= 0
*.ic v(Qout_N745)= 0
*.ic v(Qout_N746)= 0
*.ic v(Qout_N747)= 0
*.ic v(Qout_N748)= 0
*.ic v(Qout_N749)= 0
*.ic v(Qout_N750)= 0
*.ic v(Qout_N751)= 0
*.ic v(Qout_N752)= 0
*.ic v(Qout_N753)= 0
*.ic v(Qout_N754)= 0
*.ic v(Qout_N755)= 0


.control
tran 20ps 6.5e-08s

**Uncomment the following and run this spice file, if you need a waveform
**write waveform_file.raw v(clk) v(input_dec_2_) v(input_dec_1_) v(input_dec_0_)  v(output_dec_3_) v(output_dec_1_) 
*+v.xdecoder_behav_pnr.xu11.vcharge#branch 

**************************** Measuring Flip Flop output at falling edge *************************************************
meas tran ff_op_0 MAX v(Xc499_clk_opFF.iDFF_1_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_1 MAX v(Xc499_clk_opFF.iDFF_2_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_2 MAX v(Xc499_clk_opFF.iDFF_3_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_3 MAX v(Xc499_clk_opFF.iDFF_4_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_4 MAX v(Xc499_clk_opFF.iDFF_5_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_5 MAX v(Xc499_clk_opFF.iDFF_6_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_6 MAX v(Xc499_clk_opFF.iDFF_7_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_7 MAX v(Xc499_clk_opFF.iDFF_8_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_8 MAX v(Xc499_clk_opFF.iDFF_9_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_9 MAX v(Xc499_clk_opFF.iDFF_10_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_10 MAX v(Xc499_clk_opFF.iDFF_11_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_11 MAX v(Xc499_clk_opFF.iDFF_12_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_12 MAX v(Xc499_clk_opFF.iDFF_13_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_13 MAX v(Xc499_clk_opFF.iDFF_14_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_14 MAX v(Xc499_clk_opFF.iDFF_15_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_15 MAX v(Xc499_clk_opFF.iDFF_16_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_16 MAX v(Xc499_clk_opFF.iDFF_17_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_17 MAX v(Xc499_clk_opFF.iDFF_18_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_18 MAX v(Xc499_clk_opFF.iDFF_19_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_19 MAX v(Xc499_clk_opFF.iDFF_20_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_20 MAX v(Xc499_clk_opFF.iDFF_21_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_21 MAX v(Xc499_clk_opFF.iDFF_22_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_22 MAX v(Xc499_clk_opFF.iDFF_23_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_23 MAX v(Xc499_clk_opFF.iDFF_24_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_24 MAX v(Xc499_clk_opFF.iDFF_25_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_25 MAX v(Xc499_clk_opFF.iDFF_26_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_26 MAX v(Xc499_clk_opFF.iDFF_27_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_27 MAX v(Xc499_clk_opFF.iDFF_28_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_28 MAX v(Xc499_clk_opFF.iDFF_29_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_29 MAX v(Xc499_clk_opFF.iDFF_30_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_30 MAX v(Xc499_clk_opFF.iDFF_31_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_31 MAX v(Xc499_clk_opFF.iDFF_32_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_32 MAX v(Xc499_clk_opFF.iDFF_33_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_33 MAX v(Xc499_clk_opFF.iDFF_34_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_34 MAX v(Xc499_clk_opFF.iDFF_35_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_35 MAX v(Xc499_clk_opFF.iDFF_36_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_36 MAX v(Xc499_clk_opFF.iDFF_37_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_37 MAX v(Xc499_clk_opFF.iDFF_38_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_38 MAX v(Xc499_clk_opFF.iDFF_39_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_39 MAX v(Xc499_clk_opFF.iDFF_40_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_40 MAX v(Xc499_clk_opFF.iDFF_41_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_41 MAX v(Xc499_clk_opFF.DFF_1_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_42 MAX v(Xc499_clk_opFF.DFF_2_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_43 MAX v(Xc499_clk_opFF.DFF_3_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_44 MAX v(Xc499_clk_opFF.DFF_4_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_45 MAX v(Xc499_clk_opFF.DFF_5_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_46 MAX v(Xc499_clk_opFF.DFF_6_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_47 MAX v(Xc499_clk_opFF.DFF_7_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_48 MAX v(Xc499_clk_opFF.DFF_8_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_49 MAX v(Xc499_clk_opFF.DFF_9_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_50 MAX v(Xc499_clk_opFF.DFF_10_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_51 MAX v(Xc499_clk_opFF.DFF_11_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_52 MAX v(Xc499_clk_opFF.DFF_12_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_53 MAX v(Xc499_clk_opFF.DFF_13_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_54 MAX v(Xc499_clk_opFF.DFF_14_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_55 MAX v(Xc499_clk_opFF.DFF_15_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_56 MAX v(Xc499_clk_opFF.DFF_16_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_57 MAX v(Xc499_clk_opFF.DFF_17_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_58 MAX v(Xc499_clk_opFF.DFF_18_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_59 MAX v(Xc499_clk_opFF.DFF_19_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_60 MAX v(Xc499_clk_opFF.DFF_20_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_61 MAX v(Xc499_clk_opFF.DFF_21_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_62 MAX v(Xc499_clk_opFF.DFF_22_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_63 MAX v(Xc499_clk_opFF.DFF_23_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_64 MAX v(Xc499_clk_opFF.DFF_24_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_65 MAX v(Xc499_clk_opFF.DFF_25_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_66 MAX v(Xc499_clk_opFF.DFF_26_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_67 MAX v(Xc499_clk_opFF.DFF_27_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_68 MAX v(Xc499_clk_opFF.DFF_28_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_69 MAX v(Xc499_clk_opFF.DFF_29_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_70 MAX v(Xc499_clk_opFF.DFF_30_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_71 MAX v(Xc499_clk_opFF.DFF_31_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_72 MAX v(Xc499_clk_opFF.DFF_32_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_73 MAX v(Xc499_clk_opFF.oDFF_1_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_74 MAX v(Xc499_clk_opFF.oDFF_2_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_75 MAX v(Xc499_clk_opFF.oDFF_3_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_76 MAX v(Xc499_clk_opFF.oDFF_4_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_77 MAX v(Xc499_clk_opFF.oDFF_5_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_78 MAX v(Xc499_clk_opFF.oDFF_6_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_79 MAX v(Xc499_clk_opFF.oDFF_7_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_80 MAX v(Xc499_clk_opFF.oDFF_8_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_81 MAX v(Xc499_clk_opFF.oDFF_9_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_82 MAX v(Xc499_clk_opFF.oDFF_10_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_83 MAX v(Xc499_clk_opFF.oDFF_11_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_84 MAX v(Xc499_clk_opFF.oDFF_12_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_85 MAX v(Xc499_clk_opFF.oDFF_13_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_86 MAX v(Xc499_clk_opFF.oDFF_14_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_87 MAX v(Xc499_clk_opFF.oDFF_15_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_88 MAX v(Xc499_clk_opFF.oDFF_16_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_89 MAX v(Xc499_clk_opFF.oDFF_17_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_90 MAX v(Xc499_clk_opFF.oDFF_18_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_91 MAX v(Xc499_clk_opFF.oDFF_19_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_92 MAX v(Xc499_clk_opFF.oDFF_20_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_93 MAX v(Xc499_clk_opFF.oDFF_21_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_94 MAX v(Xc499_clk_opFF.oDFF_22_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_95 MAX v(Xc499_clk_opFF.oDFF_23_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_96 MAX v(Xc499_clk_opFF.oDFF_24_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_97 MAX v(Xc499_clk_opFF.oDFF_25_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_98 MAX v(Xc499_clk_opFF.oDFF_26_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_99 MAX v(Xc499_clk_opFF.oDFF_27_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_100 MAX v(Xc499_clk_opFF.oDFF_28_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_101 MAX v(Xc499_clk_opFF.oDFF_29_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_102 MAX v(Xc499_clk_opFF.oDFF_30_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_103 MAX v(Xc499_clk_opFF.oDFF_31_q_reg:Q) from=6e-08s to=6.2e-08s
meas tran ff_op_104 MAX v(Xc499_clk_opFF.oDFF_32_q_reg:Q) from=6e-08s to=6.2e-08s


***************** saving the outputs ****************
echo "$&ff_op_0" , > glitch_report_outputs_##deck_num##.csv  $$New file
echo "$&ff_op_1" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_2" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_3" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_4" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_5" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_6" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_7" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_8" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_9" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_10" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_11" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_12" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_13" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_14" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_15" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_16" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_17" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_18" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_19" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_20" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_21" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_22" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_23" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_24" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_25" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_26" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_27" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_28" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_29" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_30" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_31" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_32" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_33" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_34" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_35" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_36" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_37" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_38" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_39" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_40" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_41" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_42" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_43" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_44" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_45" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_46" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_47" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_48" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_49" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_50" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_51" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_52" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_53" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_54" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_55" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_56" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_57" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_58" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_59" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_60" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_61" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_62" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_63" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_64" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_65" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_66" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_67" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_68" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_69" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_70" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_71" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_72" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_73" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_74" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_75" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_76" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_77" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_78" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_79" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_80" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_81" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_82" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_83" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_84" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_85" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_86" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_87" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_88" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_89" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_90" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_91" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_92" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_93" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_94" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_95" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_96" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_97" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_98" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_99" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_100" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_101" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_102" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_103" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file
echo "$&ff_op_104" , >> glitch_report_outputs_##deck_num##.csv  $$Appending to the file

quit

.endc


.end

** NUMBER OF OUTPUT PINS = 105